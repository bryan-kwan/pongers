��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)��<�=�!ʢ+���#x��ȴ�jo\v�+����f�w	�GG[��m�Ce=䂓�7,�JrQE=v��dZܑ���Af�:C�M��oz�?��T6wma^bX�:ëVÙȥ��ju�[1�>)AѪ����S���L��1��`�."i�bwfа~6��D9����*�L��O�L��K-��d��22�r(�[��B_ɪ�*�����hXE�$��?p��Y�D�-�o1�x�_&���j�ˠ��u�Ù��L�#����3>\^�w}�˳�S��ev@�Y\Ņ�[9@�"��ǋ�x��sNC�CS�x��=e�*ȑ��m%��/� ,MB����P�ׁ&s��s��1�#�+Y�vɩ��[�m%�s����vN���ع"0l�6 cd''��G{V�}X;Z�u�jI��e�3[���,��7W�/%jlm�`�]�����:<mYG�0��;���2���7-���/ё9�f��oR"���X�1��w��Ӂ��0e^�q)[��؇�ջ�� na��Ep9���͞�~��K	f�v��9C��@�p�cN�v�7���K����
"<��Y��|�L�-qD-�D������uU3�Kb:�z�^n@�U�D��y����I��tz��9"���Bd�)���z��A]��N�.�4bZY�	�E]�	q�1F�Ո��蟃PuBQ��P�@���7��K�����@*��gJC�
b̨JR\����5�h=O3�&���{��>�>�;vK'�B��@M��\
�ŀ&N��\�AE�d��ϏM�E���J���/�< �Y��m�y�l�dS���Y�y�!�v����>���h+�)��耬����_�(�`ntنf��0��1��OaOƩ�������n�5bb�T�	��Qu��D�|�5��|mL"G���t*��ޑ����&�<��@A�f��*˴�������. �cs�tg)_��ן[8�Y#-AݯU��h{�W��mQ�o)A�����*{�O�(�MI\?	�,8)'KMҷ�<��U�`�p�q���b��y�Կ.`Dc����J�L^�Z"���]������\L{����\�V�TGD�]�ѷfnP���3T
��� ��
",f�l�	���9}���h������@��^����=�dx?�Op��ˮ,{g���I?t�����Ȉ�����{B��,�ǣH��߼��-�ŪrfuL��	YzS^��!#��	�m@f��]ߊ� 1Z��Ǥ�<�_��q��uT�"B��ac���[��3f@�r�w��}����L���ea�͟kգ���w_i��'��0	A�x��n��+�Զf�>ԯ��	<��?{�"C�86t��Z�\�"L:�R8[����%�H�m�	P��=ѵy���V/��܂o�J�b�,a��%�E�\�g1r/���)�*irTd�D� ����C
��������O\aq���.�O��i�8fړ�8�_b�ZY�ZW�Ě&��l�	o�]<�8D[�t��{!>�V�Ե=T��m~`�-7c2q)4�%q)���O�)4J����W�я���e1������}�FVty��G�]3a�!w��1��.-JL�l��>��V0�^�h#m�@P�~�P/m�P{��r��}`8��Ia� _��mA��(Z�?yq�V����о����P�6?�u�s-�sXd4�˨���p�Yɫɝ�7��#@�m�%$3�z��ȷ�� pa�l؉5��&F��2�(��;�t��nZ�/+�UC�.A0���=d�&�����o�˟m�C��2�-�bS,��'��h�ټNP��q�@���kiA[4�Q�\��� H}NeA�U~��c����eh]� `�Y㷜��M����E�pE_S�¤l[������݇Ȳ�F%�]x��P���5�N�:ʘ�����p���w���68�9����6'�v��v�/}���a�6v�&BND��"
˝�d����+	\�p�����=��{�dN� 	��1n7��X4��3|�4F᳄͡��˜����s�m��3CP5عP��΍X�o��C�+�B�م�D��(�\����-��N��MDL�B�g��IwhB��	�[�gf��kNf�hy����R<���hр���]�>2��`�g��N�<`/�*r�W��$�����Iv޼������9���/��fJ�^}Zh���aa��|�/I�J�4� �i��˶xÚ⟋��\���k�0����@Vn^Z�}Q��a�cm�ǋ����;.x�Zz\�N�K�@��-\n�ݾR=�z�a��>�я��j�!]fuf�,,�x�F���L�é��&���K�� 1$M�@�H�ep(�s�z|!�^hөN뿚��r~1�0��K��#���3`Z��KLB~�yA�i����*�k.m'�"
q�[�Li��q�_mJLޘ��h��.�.;;I���UQ(��m��)��.��8|��q�<����k"$�hk�yj�/�P��,%*r_��~���]2Iu:hI�!9?��t��(1��M-�_C�:$'�K]>�@�����oF�=�H��~h1�r�:I�d�Ͻ|ۖ���_�/бޑ�R�1��=g�^FN��l�����߭��k1���(%��b�b*���M�k~J�%	1k�)�X�G�]��i~�*zu��K")�,w����(��A%/Ԕ���@�ʺ�#�!v$�i��] 'I�0�4q��B��M2d��^�2	Lp?q-��c<Z�+�����NRO��0pՐ�A*F+}z���YO�y��Z��ܺ����?b䞩�D��l<3bYi�0�l����'�V��k�z���ݭ�>�Yu��}�Y���+'�
/;"B}�BB�ԕ��^
���;�dn�N`CQR9?_�?L��	�Vo�W��'��߭��$��%���>����!� �:�J�2�q	��$7�ϧ��uK���Z�(�o5�\�ei~!�� �4�'2�)�}o�*�:�����ϙ�Q�=�_Z��{۴�νr)�o��0�+�}o+�C+q=��D�=��@3���<"���WU�K�����k,�RuSG��$�iKp37V�8�=A�	���{kaO��)mZ�Uc��6a nG�͔i\y��Yʾ�,]��|M���%��A�r�&��۽� ���7�L9ٝ�b7M8�\�z�Ӄc�@�M釓�D��N&咂#�^�;���%�.?��G�1��:�9�St�US?D�	��z]y�d�2RA����"� ֖m�n���}��)�`*���eċ��̭��A��)a�z�c�>G�;��s�����24�f�,��*���Z�?ڹ@�wZ�{ɖ��n3��RP>;���mtN�e�m̀$&����������!�g6!1�k}�dJ6��ƙ%4�����P�6��,�KE�0���
��	%�|Nb��V4Y�,a�AH�T�ڽ��U����z�S~�%�]s�-1�sv"��O?zw~V�c)"��js^tvZo�[�S?�y��O�jhV(A�I� ��Z�n��u��HM�Kq�L�p�S��~N�3g��<(���Re��\�8a�ٸiX�S���g)*O�&�����rt�2�ݱ���=��}�pw���#K}l����x� �T�55_ClkvP�G�vSRp���:�'Y�nM�ĺ&Wߜ��(�
[-�)D8R�C�l�H�WiN+�JB����_M��X_\!�+�
���%Z��fƇ��II�~�w{���)f@����9��J��ip}	e�d����2��LAe�E���39�[����n��7���Y����u�����)(��W��ׇ��	c O�4skG�H0]�a����lǪ�|���@%�B��vT��I2�~5��$�B��\�YOvCI��5�ɺ-l�-O$�"9�'T�����|�֚�7E�Ic'3�e�vE�w�_���A��+���Ţzڹ����F��u���u1m�Q0r�Z��I���Y�Nc��ijh�I:}nj��<�DT!Ȉ���~�:��ջ6	��v��1��$x�ܣ����_��I�b��l��'g{���L�zF0
���@���qT��e�C]Q���w���j Y�����Q�O:sc�\��Q�I͜�?ad�43%�U*޴��hҨQR�]�z�ڐȖzX�[��Ԕ��#H�&�D��u���,)!ĸ�5|\���(�7w�Ij�X&��JS.���� �Pj|�e���to��k�0:g͑���*&l�=�z��-�)ם뗀��@- <��q1Dx�<�+�z9�y�0����k,�Y���>i��i��XPY��aP\�.�m]�*��X��q�Q�B{�]��K``�^�UT�;��\'�K����])���m����/��\���"�UQ\���b�*�̃��8�}��W5�n�:Pj}>Sn�>^��We33��O[��Y�GN��^��ݿ������H^���7�8�>΃�37i�����b��d��P���B�#4�TO@L�B��T�K�B5�Ew��K��eC�;���T�������l4P�Y�:}� ;�3��;���+��ɽE��2 �$֥>�C_��?m&��o�n����'!�����x���Š7����o��� g��l"�
�P<���J�TDs��r�'�>9x)�ꍳ�А�\�ξ��8f���KS�Y�ta����[��5 f
֕��c��+�@���R����yM{��S�-�V��u�����Ǚr�
����얚4��	^�s��z�=���8�6*�I�p�s�
�����,R4䵦m���X�0B�����*�_�l����	�����`M)�6��	e�s@]��;�@���4p)�;��g�����D��2�>�{F�9E��y]&����\�L�����3ƻ��:�2Q-bc��1&͎>�B�� X�d�����F�7�4���Q5��9Twd#�F�tY��T�sʼ�N�".���l��,�tu\́��Di�cAధ��#���_l�#W�7x�0N�(��� tT�������d���l]|o�dA�fQyb��X�*@]V���w����r���|���������T.��� e���-,����I��3��^ �6dȖm�e����Ȩ�-����&�{�Χ�wW�S|V,�j�c|ޞB��H�ar�d�����2��~�0J�9� G�s*$h�o���~ae#�y��^ʒ���{�t=�6��d	~���f����"
��O��巊|��f�@�*O�@��_�����֖t�����oA�R���JNd��PR���s�)�^�Au�#
��������>�M�L@�x�	�w�w������!B�"�`[�'%��e�S��f�zQ���*/ɛ*�)k�[�<��H=]�IP��g���w͸�w��z�N�i��u�)qO���Le�ߜ�9d�� :��������]����禽�aG��i�h�
-���B���Hi��4fC�tM�b=�
gK��C��p��"dM[��n���~9eo�?��R8A�#�2:*�r�-��K�t�&�����y9w���;+�.$�Tvcb����ڻ�UqL�E�v�+���%��_�1O"�Rƽ	�V�l�R��$��cL*tA�������\���+�H_�s�v��k�`7RF��Fm�9��4���ө89m��,���JI�e�P���*k�k��E�{n���`xi�t�{�:�g��a6�+%���r�{�(l1? �( XB8t\횩��&��1:j-�j��Ҋ"D���qH�e}���A: ����b9D߅��^����X	���]6�~��3�4�8:L��x{��2�jc�q��	�<�s֠~�i����o��[L�uȾ�k��m7�^�|W��8<E����u}\��3�@�'�=H3���a<(���~0|�2���Z�nv��0�Ar�T>6h�p��^�)�%qhK{v�'�[����;��ͬg��v���B>��^��������EfG�FR8Bڕ��%{����y��\4v�ʕ�D#(��_�@z;�p��>�֬�m�#,���ˏLL��9Q[*�:ڀ	�����LZ8�-˕��˻^�KK�� -H ���A��xr�Ef������
��h�<�n�rq}������B��K���Ӑ)�: f�������B��4�Wĸə{s�gH���B��Vy��rϷ���F��7�@n+����_!}-|�|��n�]s]1�vRi8�m��;�:/�H��)�g��F��k��	o�����v��r;ei_Mp朜�f���?���aj��C�at}��u�/����P�-���
^y	U,��v�s�E��M�r=�]MV��&c����*!�Ez�3>J(�5l[ѥ�
��j�M��Sߚa�8j��on7� ������=D"�1�$���s:�*��GAr�-.:���)����%i`�+y)���M�/������y����dܾ�4�az|�5q����\W�$�=�LJ�6>*堥F`���+�iy���o
��Q�S84��_�4.�#pG��з$r�oB"lH�MD���f��41v,][c�磟�]$^o����)#��<�ӳ,C6���Z2q�mc�g�,�&4f���E*D�������+qA/(���	�P�q��Ц
ځ���3�V�;��em,H�p>�h�m������AbU:�]+������N��Bl�Tgyz5�F�����V�hk�u^��^��`Y�1S�U��Wc�6匑=H�m�kL���[e�Z�7�����ga-��C���~!0��7�1K�M#x�L6t��I����^�*C��l�ʻ���7�1���{�-2�j �m�w<��7;�̾��]�ظ�Hx�F�8�r}�����^8K���+@E�hM�\NE�F��'�ԌضzsHק$��^#�2�߯�^�rx�?�L����J���6���F�Q����Ti�sc�Z�&k�SWS���_#D�69ʌ�+�z%����U�� ��@�}ɲ��8�?v�=�4�V3��@��j��qY�N���,ҟ�wʅ���Z�Ђu�� �n�eOY�����r�#��Z���~���G�x�S��p������,� 8�$�\�n��q��ɢ���:��D��߮%4+�f��>��C�.���=@ǐ1�oH���&
+�ѳ7]*^\���Y�?>�rB�k�r�b� �_�qH�|Dli��ݡ�������]F��)�ĿF�sv�!	ǫ�a頷'+�
��s��a�Pf��Pe��?��K��$���{N�*���}gCwԃ�p��q'�袝�od�tU�?P�ô��k=d��=����.����z���m�����\�2��ж��6;�F}���u�(���K��ڑYé���	�"ף�O�T��4����zr	EV>5�Y�Ovd3nE�ň�	`���r�C�\\���H;>K��v;��ʄ�9�-�%B9���S��]B�2H�c64;Ѿ0w�B�.�?��SJf��INR���� *w�J��VL�9�����`;A�2J�O��h��l�͢B9{G|E�r�P��7$��B�2L��z�_�Z�u�T{z0f୔�jO$`����PE�b�1%Գ�h��(�2�<:�g�e{;����=�g��)��C�D�`�0�3!�~0fB�̾�d1���6���@�xyr�/~ˡ� H( ��5�}�8������cЋyzڋ����sPPP��&4j���a�W׫ gR2\"�xG���7ج�"3�#*��-�����Tb8�g����|a*+���C�"�{H		z�S"�"{vj��o�Y%1�gRt���_D�/M�B�DA�B����I`���<��'�R� &	.�~���9��d����Z��R:	m�ն��4����
���8��8�H%�����5ֆP�mNt)�b~�6�~���,$��KT:Yک��9c·���SȻb�ű�-��Qi&�]���2�$��ڵ��އ>p:�2�0���?�������2������,���R�!!�:Ȯ�N���9j4�t�Χe���J>����Xs�
�+���z��nE&K�Z�
��ԝ5��~qF�ɁV����mWw]�$�V#�n��L��Gz����������m�/��	�WN��� dG[��r�U? �ns�\�G��M�vz1K6G�������y��r��$���o�=OI�A>�!�p�w��/��+7A���*��1$����RѶ�_��7T�Gx�4f�oZǪ�Qu���V-�VA ���$C����H���X��[*�j}w�6U�p��.�U�Y�ꉃ0����r���ٽ(pY􇜋���m	T���"Mh�*f�����B�+ܖls��;�8�!�	� �-���Kj��8�B[��S�#<љ*��4�.�OƁ����6��d�(�J�W)���CF�h<�9C���!�;��Q�
�������|��V�7�H�pD���(��(!�S�� ��J	7m���ܾ�7@�mV��4���!�Юޅ�;��!��g�% V��Y���0�vg���i���ow��\��YsFW�o�w4����9��Ф}"F"��4x�b�����ܿ���~DV�b����k�m��1���87۾B[�J���(�9+�N�a�d^�S������n�>�8�I�;�o������ڎi�}D2��¯4�HY���ܟ�C�ƞ���D".�<���\�p.<�ך�V[�$;�Y�T>����	1����0{�m��V�9gP�|ɠ	򔔷^��`�����6�ŧ�e��Â1����O.�$�@�<é"#>�ɨ��5� IT���D���R��҂$��O����� -ၙ ��0�:L�>���u���U�_F��``'�Q��[��.�b�i�R�	�f�i���˶#�>y��#��s�����z��&��x���tx~8�Ķ /YU~��������5?rU�U"���'8c�2�fT��Y�bk�zb�职�J��{Վ�k�/M����a޹2jflW�eRS`EV(B��_�8iU���h:އ���h�E7#���RK&��L�ރ'��ƒ�=�<�Z���h=>*�lF��k��1 �!�8��X�a�4��o��ϡ�\�P���Q�w�oD�R�14Վ�ػg߶w��ލߢ�ַ`P�<s�p�#����J�
��߶�#�vxu���~u��uO��y�S�N�D���Lk�s6��`|���0��*���3�׀���ws����wԶ�����]��.#�,��Տm0������I�̇��@#i�eA�ԥ�QE�v�c�n{�O�²�b6����F�V��S%��:�ce�K79I�p��kx�W�,(׃��V�}oɿu:�+�Fh��&��>`����o)��_.f�DKƽ�(4��`j�E��7j )��*� �9���{j��xʉu}��y��hu���ĭ����t5����4�^�D���@tye㝓���ą::D��j�U0
ks�L5���9,^��-E�'b�:��
�ȗ��+�}��β��9�6��T��y�p��� ��p���tAܖ��s�zbq��}����F��}���6�H��㤾M��rb;�a��'db:���b��t�0A���b[��xGH<�X	�� 7}�N��-�x��
�ŷ�Qy$R���H1��@K��))B��.����;A+���͘��G��O��T�a:��cB�~��=X���v+���7�j/уn�{��� 77�m*X+qG�1��m������]��9[P�mܔvB������+���E[�~���D�ȶ�b�ro �Ǫ�g&�<p���d��'�j��C�$���4#��_��AX��^�u!_ YŮt�ɏ���3[��f^�Gg��~������}�-��q�[ �\S��Z������ �n_f�ױ�'voaK)p�q���q즋m?�2�"�i��~(��8	�=- 7ܓ�Q���lcp�q)�K�M!ɴlM�FUΓ'��6��ɕ���/�+&����|]�i�9�>��mC�5��vO,#����r���k>W���8gI'RJ���ٔ�������'n�q|�= eXY�&�]*{��@e�����񝦌����d���U�^+=yͨ���2	x�W�]0�3�o�˃���� ׀���h�!n��3)D�
�v���Z�V�b��Ww���u��dn�&<*/�z!&aAl^�S|�(��d�4l�V�b=p=Y�Z�'W���:!w^�/������GX4����|���j�ui��*P�5
�4�l����ںR�g(���
ɖ�Nrw�P��7������Ʉ��ɧ������f�'q(PRŧ����c�y��@9XFLA�����Z��ǉ3R�A=p�}mU�aAp�hQa���}GT�
9�S/Y�Xb}��w��(�LTcX��!��X�)�3��[&�l� /�o:n�#Ue4�_7��h��2a�3�t�2 �t��;!�*�������*�E=ύ�d��v��Q���e�6]E�u�����ar�Β����;��j�Td�|�B�0����w���r��	ض��y��/H���S��W�EV��4��q�`5�wP�r�Ԣ�^��7�����V�V�)`p���lֽ�!�6��_�^�4��z����T��|��(auϖ��$���sr�C�̥�TC���9蠑�S`��[�!��2���o����WؤǌL�e]�k8t�H؉|%��!�w`��`&+�`��pC��<<���)��,��Q��]l��Kz��4��������!�q�G�ͤ�nتS0a=� \[疇��h���p`;_��	�]v��,D�X.���%eV�/f�0���T�2��N���	ً��]�؛�s\D�DdEb��C�b"��ٺx(-��$��9��js}Ǆ5�$h¦mBU���Nr�Kv��r���g�Ά�L@0sDʣ�Ƞx���C�b�Z�6@$*��� �I
���o�y�f�L���,�X��H<a� *`ɂ? �.�̄>b���O��h:$o��� ����z�&CfrP"i;�n�/��D�l���P� ��
����j⥈J�76}f�n'oP�b���)1��9�
� ���y��b�Ė���Ҽ�~�eK�m?����Ӟ��f���%�8\�Dp3}�1��o�@�f���s��$�^�E�:���
�C9g������-�﬋u��}g��
QG����AQG�5
�,��-���nt6� y��H��oJ�V5����8�ץ���og
����Q3�7Zw~>?p'���(�-ߑ��F�>@�#��{N6�4��I��:����[�w4�#Ve��J�HC>h�/fցg/������2�/>j)u�e�Q$;v�#Lv���l�N����0֗\�7�Ҁi];G@�~��!��݌
��Q��;����	Z"�.����J8W>m<�ٌ�A�B�tz�*���6����:P�����3�����J{��x$Tt�]�u<A��,�[���`d�G���ps�7*ָI$�����Cu�9Ea��� w��ov˙���h�~��u�<L�� �}����jbAʷ���C��o.�k���3 �K?T����˚��֨�9,���L/1D]�O�,�ځd =i��SȐ��:&á��;
�s^���E"���n"���Mz�nE����2	Ai׌ ���:�^�i��\���?r�)��`��Ѱm b�?�K".�5R�2Ŵ���=\��o1r2��p�D��-��&� ٽj�>�.O	j�D�Z�W8MagEA�B���,�ݷ+v���JC�2AI<{r��8A]L�w8�P}��O+���so��G��<?�`�����E�`�=;
���^�{MpFE]|e�8b$Hj��Sc��A	�'���B�勤�"��e�#P�Ft�if�Q!Њp�6?�����y4Ĳ��^4 N�������i���#�bv�u���=4_lYt�;Z}t�z	w~v�T�P�h�<�K-����?ժ���[�k2H趂CL�_EZQU�����o9,3w.����8soc$�,:Π��9{�!�m�� &i�;�E`�}�ϣ���P��I�v������(}�	 ��|!�-$Z~��*6�E"�dߵ�۽H(��b�+e���}��I���+�w0�'̼����I~h�K�0�!�[GJ���2���ą'e��kX�o9�m����{W@�a�����=&�֌ �}�W���A1��E�`L�ȩn�#��Q9�e}����_t��c�ä?�S��د�d�3�-�?�p�²s4����*�Du�ۼk�DJ)�ɮ6���S=1��7�ߗ����G]�>���@4��ɞm���OBRe�y$6�---uJ$I��O,�eѬ��O�l�YDZ+�C.Irt*U��@֩����W��8�#��M�������K5��f7b)�d9��23[]�d��)�Y�fF��H��N���٤����{��6烎U<ᣝG��MY-�p1�]Ӿ��'y��)/�E����+G�6����� �e��w�S`�N�=�v2=aOu]�6gO;��[�1�F��2��o��͎ �&!2Z�8�}H�au�L�;���ź��efo�W����d��2;�^��vE����sD�!@Q�@R���������(��R�=m�I�+����3��Vu/8I.A}3���3C��&vo[b�(��H�� l�KP��p��$����)+���$��&D�U�G ��H������F��c,˿�����A�IY.��
|ba(u��	]����p���N*KM��<��1��~شm�r����!�P3,����Uo�&i�T�S ����٭��aR��֥��5��][��������kx�Y�����H>��q�D��%U(n��1���@�{���t��j��k�tM���:Gu1�lH8l�&B���B���{V�V�Ys��?�սFTe�)M;M�؜Vc���"eq{�%H*���F���$�؀�����}��1)\���;
j�F�_��*�8��۸aNεx��;��/�G�MP�R��v	r9Y�u�gƑ�X�s���`����fD�{���G�,W
�D%_�����W���G�CmF]���������.�5�K�7�=D��;��HW5����[#�C��3#�;u���/�[C���\�Mm"xW^�dQ�����F-��w̖��-�bk\w䮸�}��"O3��D����Ԩ	>�(�R�U3���0� .�H�$`q[������e�:����L.��eX8�C}H��]��H<s�)+�;_>��O��cG}}��|��%LD��,$�&��Jgvg�sD��D��ol���оk�~-z�3���6!�g��?!��@�u���yϕ�_|�r��UA��W�*��^�G�?�K�� �|�`W��2?_[,2�Cu`3��=fe��jh�8��;�W��GfMᬦ�MT���!T�P-l7;Hy�.�YX&oog2�R�	�:�p�����?	3;u�7�,���W�p.���;�]m����5,xy�pY�DkY�"t~��#f�X3�+Uu=Һqx��⇕'��c�C#̈�U˂<���}/�(f��[����QN�8�.7�P��� &�5ω��
��^����Ab[���0�褓���AUѶ��GF�&UT̡�0���:G�n���"`�����6��HV��rbZ�h7�����S�__�ۃ�6�k�牋�/�g���*s�����P؛�u��g�2�甘q����VȦ��Ն�����)��Y����ь]�b��3�ݝv����¤����c-��ٍ��^�47q�)�GXE�4:$����ʶ-	�YĒ$�%1_Ș�3��XTv���Q���ާ�	�I��4�͆ž�+���}M�6�uZ�0>��t�V���Pf̟�^�^���N^^��9G�dt {P:H,�CpYϔ�.�YGn��Å�3�wj�䓗pIA��Q��3�''�J ���&��T���
R �8s�[Ǝ�='-��޷H/P1�RB�O��o�����yv��{2��1�6���<�y��k�e��!!*�8ԙiE+��;���n=����t��y�%�Ȃ���a�V�h�'���R�[)�oi0v^ٕ���m�M;��٤1��]�q�u\-�x�Z97��\^CEu�S�wŔ1Д�#|�z�V�6@m��w;�e��J��a1��g�+4½�h�~�"�e(F�y��{�3;�t�q�@O5�����?�[����_���x0����^�"�`y�p�$L�$͉��� ����*�ď��&Q��^@�e�vK��mq��0zI�F?�n������'��A+|	:��6�C6�oB��dna�p��	�6G�^vV�;��	�z>J~�F1���VM3�`��
l\ku�'�����5;yEW����I��M\��mn3�Ef��C�Q���$`�<���_�@������-&@��޿�/�-���\�!y�,oN�\#���ʨ�榊�9U�,� ����O%-_.�΍��X��x�����x+�!�u:#D# �րxxY�S:�x���zzq��n��)/)I��g��j�I\�%t�A�	��Y�wE@L��J:��Pd�m���6�&ˋ��ʪc(.����¡��γ�&]�W�O��|���OP���ڨ���p��{��Ls��v�60�x4�Wh�]��1��2ī�]�x����S�ׯ`p�p�L[*�r�lF�+͎X��Dh��*:L����f��9�����0i����r�5��k㑶g����'�Q|O$[A���_w��4�	�Y�
]좎����	7A`�
�F���u�v�u�F���y���;�x�9voۇU12@�.v@恫�V��{�wL�tڧ��p2��K�n�*9W�] �n`J=7cǌy�t�
� җ6G������xw]?�O�t`zⴡ��ue=�c6MFx�J�В/�{L�CVDBi�m̠M���Z�<��21dM 凨�"_B� l�X�k�S߅�D��1C��J��mԡ��h���Ѯ�Ei�O��(�.���*�nV�H�¯ ��QQ�(@��.��<@�lwh�:�v�>�vpX�����%<�_�:�T1Ƚ-�e�Z��4��:�'�%Lc��,���00z��.��i�����@ݢ[׮6m��xl6^�K�d9ӯu4f��oz�U%h5����ܓ��H|�.�QN<�ĥK���l����Z<����t�R6�m��@ŏrg&x�&����'��h��R��[J %�����("�9�5�+��v�nITd��q7[�Žz�FB����1?�@қ��c21���R�+��R�f��tE���E���dy[���S�Z��O�#Y����A�Q���3J�T�N�}(V@Qq?纤S=����P{0
We�_G��z���{�y�U��L܂fk�KJ龪j$F{LKJԐ{���ɮ
���7X.��b;��8������ŭee�3����ƞbuj�mQRd��Y��wKà�UT����_@0ݭ6B�]c�~��S� �PS.��^��<9-�0����0�~�.�V���!��j?̕Eo�3aF��<��8!W���%���s��,�����Y�_wX��C���6�~���L�u_�4�!xʪ��o�ؑ	�c�N2ї�胳A[C��. ��8u�8GM�@i+)�϶��m���+X��3���f�+��&��0_�����6Yge�{"B����P���3����y��&��ΊF��u۟*�ţ6��ͮ�+��n�ֿ9�i�߿8�-�iI���c�_F'*���F�6�:iVͪy��Ȥ����&;�i(-�f�7��)��5���Xüt������o��C2������-��E7i�����L�\B��Q���L��|k�iԺ�17�">�ab���eW�dk���[�P_����5GS:8Շ���*X6T+e G�Z�V��~��r�=�5@��5�7��}���O2�9o����c�A�4� ��V�7�>�{������4��m��H��̨����2�71c�{����@� z����������k?��R-D¯v8N��kH�]8�+��$��B_⿝1�i�J��2Ve(����(
8_�o���I�R�K�`|:���)�2O�o_*����`6,L0�Cҁ�`�J:����mj�W�5�"�Фb��@�F��'�y�ؙ��kI��Uk�@;Y���Y��I��"�O
���	�U��谡���!� -���A!��st���:�=�FP�+��W�J�q��[+����jO�U��?�<��