��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)�2������2p|�t����:8��P�_ ��U��bkS��p8|"-Q�>2!��l���z�NG}���V�L��j�B��t[���'t�m��j��=��:��M�J.0-�+���0Y����*2�y�C��/��l%��$E�a��N>��>�;\�J��4Hh��X���U�����S�(��_���:>���DƩ����-AU-��V�O3���'/�%�:MQ�qͳ Z*�&�'�^�BT[ ��{1"g3�m1ă �=,�����W��f��T
],�s#.ϧ�F��]1���&5� �#�xk��O�c.�
�����N!�MG��gہ�����܌��%o0�����4��Y�Sҏ֎$I0���<����-�yQ�}uYʨ�ԭ��z�>��N�i���x;5�� ��w�5f�fЕu��ɕ�}Bf�3; ��FE~��o-!� j�����Pn�9O����;�o���򈤣��xJ��ܷ#t���� _8�#�ql��>j�y�:�;2�.���U�����'�=/���=*��G*_{|"�]���.O	U�j�=�h]���}pV�J�Лd�O�����!�P��q�=0aw�ͤN �,Y9��w��*����F����>�/��X��G�W{#0�g���q^e�K&O�[��s���{a'�����S��׷3�zșc�zM��"�o-����~]�[PQ���ۑ�(�#�2/��f@�B�sk[�W�]�yt����L��×�EQ���p�n�hΪA�,ȕ��m���af���cPl{�g��"Ԉ.��c�Wnl��W������//~N�.�����i�ύL?�c*&O�2��%�hn���ʞ���Ѱ�-HMB�Eb�JǊ�q������jn.���fa/�y����P�JT�}�ş�M�4~��W��@�y�ԭ;��=�xR�S��o[Sɭ��}��8u������w?܌Ma|�?��#r1�'��C��_E-�P>���AnUHB)�7�~/I�1l�[5��Ə������.�;�(U���)�wҜ?۳F\m����E��(V8��-�5�<9����P,�1�'&�ș�_�ߵ������/����!<�Z��z�~���Z�`$Sm'r��۳Z~��$��a��N������B�n&R=E�|�����^
��UTK1")�[e�7�.�(䝋��qFn���Ut� ����$.�$��HF���2�4�C�g�7d�0�b���SY����}h��2�4��q�r��o����F��'��I6�yUMM�x �;��fz��}��׭��&�jl:���ѵm����c{�maV�º�j�x�.��k]���p+�3�yd�@5��:�$�㥋����C�	^�m.��`�� ]�?2'��HE�QH�ta�8p��#IQ(� �g�Gi�4*��M;)r����N\q-3�\����h��"W+aގ�o�]��R��O� �"g�T o	,Y�R]=5F7ti�L?l��l�kی�ZQ�Iʕ�c�_+J�=���Ql�7�s�w���UGͣ6��f*��:]���rl�D췜pɖ�KM�8l�mj�}�Z/r�\�Y���:�w�&	Lp$d��E�m6��]vjra�2�M�f���k���%���űmؘ��J=W�_ͬ��og.&9 ��Z2���������>+E�X�܏+��	�=)��iz�6�Z!�T�g��+�����s�o@QJH�7M:R̤ &z����5�@v_j��u���{V��7ޚe���]�����q!��ui4c��Xu�.��m��X��K56�Q(dgP]Խ���[�� ��SPj\7v8b*� ����;��9Ɣn5
h���$SB�߹�(�"�I�I����g��{��_ʽN{�'a��L֙+��>z)dD��lxY�A��»�dB*�0ȐZ�#%�M*"�e3Pw(�|b>$���k���y[ $�����9nT��\�R���z�'��$h/�E����1��L�fۆ�f��k*�SJ>����Gh�9�IS�Nઝb�%��怆_S�	�*ہ�<�'*��H;��i���);�a�M�!U�R�|���U�~y�e� ���Z����� �
dp��Oms�]*b�<Sz�$���W- �DTA������R��oo����|�`SO"���y��ϭ��U}�Y���q��2�� :�[)O<)Th3��E�~5�R�}c�i�Լ�4ƌ.�#�i_8�x�T�u���'BtEsIw�ى��S3w4���>��X���k��8S�����~	�g�kzE% �L�Hj�>-t�HC'���s��o�8��m���Q�H9�p�?�0���r@n?h��a���Ҫ�;�>����{��e��q5��4�㗾Z|����j�u���M.
ԥ��A��{��M3���m�_�ۮ�8`��� ;A�I��1�X�YU`�;XG�O\)��}m�����B��8�~a�0�{9��A,���!A�[�j
ϝC��j�U�PVSJ�0&��!D넛F����kS0U�覨�]纺E���=Ǩ��	�PpF9qu�R�����C���l6s�4�zV����`~��y�L	(�Vf3q�A�A�{��ؖ+����d��?��R���6�+�v�ܥ)�f����I�e�j�Ů5���/X���8K��Jں����jfvu�h4��j<9���d*�H��B�0V������?1&ε��?X%R���%�f����z�8�%��&*�2����H�w�F_;S\�cXW.��L�X��ls�߈�F;,�'�|m~�y�rR�6z��yZ�hDh��ֲ�?C�	3q..�ܦ-wP�X��`�q7�P� ����_��&n=-��yy����<�`q�\���+o����̅�h�q�LӰ��꒫_~qǨ�p~��aKg2�J�ӕR�vb/�� ��6-:6Ҧӧ�U/�O|�0.b��+�M]�lX_pE�	��a4��)���YM��?��|Ԏ���[�������@~�����+M��7L����!8��	AW>l��~��d4�M9ꪐ��cK[V}ܭc,C�6�C�I(�����D-/.����,���)Yi�N�����"�0�C�uk{������U�q[Q��r�'����b���O@]����N
8�5�di�C�)�Lr���ψ��:�G��Õ�q:;*.g1�=�oͱ�ղtIh�v4�/�4�ً�<@Jo{D�כd�G��	�&�,j��O�0��v���F�)	������ �l�M�w��N�Pf�%�̶�B���>.��ݻ��TGe�?�|-K8	@�(��)��n�[C�Rs�h��f��>t>?�������Ư�fdUm�ʻ3�W�/�~ET
+XO�3��%��֧� �%��մ�NL��E��Y�;�s�� &��,�.���d�$w՞�x�[��>]=w�c$U�Z����݉
��#p�F�Q^����g/&=/�C���D����K[�G��)��
/x�H�Fb�����	Mg������_*�7�[�v�9�����T��l�3�١�N�ǳ�i����u�w������M����.�VS���7Y��j��=ֵ�͙N�G�s�p��8��9 ��~�g�!#LdC�Vj/�	Rx3�U�^+0)��l��,�Z(ӫ���e����
TŒ�д,���Įt�#'Щ��N�<��cf�V�F_]I%H��8(��u�!�j�/nfެ��9�2����F��N����ͫd&�����}��*�n���\rB�� �4	�&�E$2멊��q<0Z�C�i$~���C�7��+"�Ų��$;��%z�7U��i�D�5u���O��ް�}>Jg@N�O>;���W��Q0,������ƞ��Z��m6})���ҋ��9�c��h�J�Dv�>}�aR�s`Iu��/6��Q���~��y@��)┬�j	�q��\�`Q��=B�38N�.�r��,���m�|/Ҕ\��(0���8{`wӭ�Y �;8��.����{1�N~e"���
��ǣ��Y0/	�� /���~����­��CHԄc�qǙ����\Z��/7E����$W�edu�˖��q��\�Ҁ�$�b��2��~E�6�6h(޽0GWA5<�Jzn����$�2"��Y�+����EwG!�)��!!��}���6���'HY����ZT^2��:N����\���2�!+m6U鸷_�=�0U� �C���N�n<�o�����;5^��,|�qJ�U<�\����yV�����k@�?�"8VL�8�N�{�&� �}�⒔���
@��:����S|gH����흞�,͟O����6�I�[=��hK\4�mϘ�C����'v��v�/���r�`��	���%B����!���u��	��w4�'���2�D�W⁽lo�W�?��|�\鋅��'��-7Y������2��|���D�"��݅Z��� 1f��?�s���ŵ=K�М������y�kl7������b�
�!�>P��HV��"IMч��:(MwW��L�cί����(��/ZR[:F����+	J�8�\����� \Z�� B\}���r�A��@����N�*�Q���j����1�l��n�HKГ�C2,������*,�et1#�N<H�窃`���a���;�����T@�3��Y�$'C u�K4�Z(�
�t\B]|����o1�N�w-��̤�>�%w���_�I��w&���S�?-��J��T�P;N~Ǿ�褻�p[0Zn$�n�P O ��'֏%��ybh~�t~;~��x��r�������Q5��+�Z�À��f ,g?;�~H��s�ӖN��:�e���"}z"���qj����ְ���>���i	GqڦŪ�4��5��؜Ȑ�:�0=�w�� �+M悔���A *���V���3�3|����	���y��z'��{-х�7Xy�GMl�6A��qnc��{T��������Q�(A|�����{�^ϧ��M�Z����_1�Yh7��	�%�o��2��^F�NMu�#���jg6�U�T���Q�.)�x_l��u�	S����&��{[A�#]̚y��p��V�npU�֏���l���i�����#���OH���FwN���o���O�v�b��������^?|{��5gKSCs�c^&�U��v4��:c�	�R�����=u��8s�IQa�[����G��g���x��EtvY���3|���6��|�A��k�+[���8	�����p8��ߠ6�3n�]qZ["0-,����^��a9_���h���lC�8�Y��MFjT�.t�EN=��'1Ҧ�$�j����"}�G|���l�������N�.���R=�ƛ�*_�����3 |�(�ĕ��d�W>�{�Qy��P0����?X����