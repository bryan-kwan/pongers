��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)�2������2p|�t����22���TO��K9��c�"A��{,,�BF,8,�.4~�n�a}��B0E��W�Y� ����Z'�2��;<�S��3y�}��SSi�*g���T��p��{�#��	�hF�K_u"��Ir���&Ŵ���ls�n��F����4]ɉ����СM�ˎ0�g0r:u�f| ��ѽgNX4�ۡ���,�K��^nXV�]�u_�"x��<�^;m3��w6N����x�##��G�U���x�a�j�L�6q�nC�1�&�Ӎө�`�59�&�|=��85R�$H�^]汁,��V�X�Q�˙.�yN�fh34�/��N��;_9���^|\�~�^�z&�=YI�e�<����U��8�q~�SI�T�	�L�L@!�n$Ʈӑ����%�z��R�+���?�:1�Tp5a�.�Ɖ#ٺ�o�́'��Akr{��y���� ��R	L��XM4���n�ж���H<�����H�D����&m%�ضs�A��%6=�Ҽ���4��||$po�&
���O���/ S�Sb�'D��<��U�sW�
ҟ3���tl��������QW|�'��;z���cIB{6�^i��n���x��$�SA��Xm�����R�T��I��������}�E{�3e%��|�Ňk�..��d�14.Ф,��RC��*.�8?�����՜;=���$�����R�����������q�Ȓ��7j'4>��UZZc��|�R�P(TY��.aoY���\��C�By1��_P�e�u�k�i����=>�)�<�G�3�n��%U*z���_��F��|4����9f�]�<S<����aK�5B��D����T��_��4!��Ｏ,ڦ�$�:��b!�H�o��Rh�#���!���0�3��(�LK��лLA����:���&RCp鈽vc���%��w �T�$� �"o2�����՛���nj���7	=��@~%s��!7�ٳ�^Bw��g�SY�������rv����Bt#��8Ȋt3�^mWU��h,��|呅���>ܶ��Ԕx����ɔ�#]��@�6��:�Z�x{�j���K}�*~�	��j���]c���Q���r"$���_��g�"�\H�$)2e^qmq^A#:r.��9��z�$5fX����ϕ������ժ�e�O}����+޶OZ�[my�C�g:&��k�_�iGK�݁m�(�VF��ʍ�b�0MY����>0���9�SfY�����&���IA���&���������I>�����ս=ԁ@���aJ����,7~��W}4�5���������`���^K��,��k�M3��w$���
Ǚ�eBA#�k��h�cD�&]~��Ĩ]Ϣ(2[��Lk�ޑ��e��7�A���ep�)&�m��������_bG:w���`��b�Ƣ��=<r��
S	*�/�4��FV�s
��4�^F��q�v�o�!,�#�Y'�T�F����ﵻNQԧ��T�U����x�\��� ��m\�'���zt^R��64m�;�@�w�C��8[��J8��TT/���w�rS�6Y�3x�5��W�����F�e�&���
$/1}Sݙ�;}���p�"4�QÛ~A��}��tW&>N}��I��Ĥ3C�\����ٝ�h�H�������휲p��Vqu�Zzj��]Ēw�Zϭ�O�ζ�8B�����n:�?�v\�sA������l�Q5u�+�N�@}?]�9�$���_����+Fv:`2�Ҍz���H,18��Z��:�gΰ�'��wn*���aҺ����u�W/�uZf�L��0�kU��kO��9ԓ�x�l���h�����M��<8��B�{�lT�7ņ����0���C�5^0A�
���"5�;!<��Ok�v᪖�ѹ?L�NB¼Y��;{�Q\TI�ś�ܛ��%�]M��n��ᤥ"�$����#��,�軹��_b��c�K!��>�"i���蔾�p_����	�{�2�>�;�Q�I<6�"���ʯmZp�|�j-iC�P�W�!�j3Ⱥ�R0/8^d�_P�n���q2�|rC)���\m�����<�f*br��b�� w�zˤ|$�a0��bh���N�#"���:f/+w�%M�J!�nW�CD;�%��#<,0}������>*��:1�X?���PQ�)O���߻�X��/�ct��h.T�����;�����&S����v,���X�4$]���ö�B/��>�	��w�5L��A�����@��l��N��
4��n�h5���o��т�Q�xq�`��
�=������'���{X����/}͸�Er>�{�ϑ�<~�'��	���KA��kVT�UJ������`��'v�:����,29����F�عbB���犘?�����d�a�9�q��܌��cÛ���!��O�
�G�㓺]�튑�?S�ӓH?�q���:C��b-_jI�M�=��~�B�}�>��Y���Z"s'a�s�j�U�++jbl��ʚ|�� �A	�P=wIl��4�3r���b�2�f.���1{�`8f�z;�!���
kB��蕨p�R�%$'�Us�d'�I�m4�z$���# z#�O����QW��c�"杬f8v@�N<�a�n�ih�_��(�	�4I�k!X�+�m��x[��� �4���t��=,�K���7&О� ��4�@����C&��r���E��������ᣦ؁	|�ó H��uo�{j��w9+��#���A�D
��DF:���1.��2�3���v&4��|BuU3�h>�_��3�v4Q8|�Bt��,�Q{T����'�x�P�<$���2u榚H�9U�:Iw3���f���Qo3�1ǐ�UF!���g�Q�r��?%�$�)�����i2��rD�Ѭ{�ZiDab��8�	��H����+i�ݡ"�<�#gn;%^�V���[��U����BH��'��\�\���+���n,�m6gv��8�!2���fh�;�RRm_!ȿ�/]x����1o�b���j*����s}�S, FW������x�V_����|l4�!`���_�g�
5=�L�b!���[�1�Gw'�:���v����ן9��<�3��gpN��l�D�A�V��X\��Xލ4�!DY�u|c�k+��D���{��Z��{l��|��l;h���To0!����+C\tͷ�(����hkV-��-�{߲D����.#R��t�wƝ������u�϶Yc�Y<ͪ��U� �Y�Y9�l>A�΀���B�߈б��f=�	�J6�l� Cs;��}�ڨ'�����$?{�W��?تw\>�_�f1�����n��ѫ��n{n�C,��7�$�濘K}�n��<uʹ;8wg`�4V�m�	o�VޥSϰ�P��V�����r];��h0����;��,�Ia�(g^�;f&�DҐ��� #Ȇ-�h�j��������I�T���2,u5g�T'2����FJ�@���9S��fe/m=�����7!��=�D�>�D����� +��RU�Z32"w
��X��Q�՟7Ŭ_f��MAMH��3�~c� �*APgF�t/�G�T�?�8�{�ۯtVeV3b����.(7����1�Zb�Q #I�[�M�8E���� %�W�9S����)alB㉄�tR��.���.���xx�-�!R�`T�eɱ�f�ט�rȏ�*|�e�[�	�n1NW�D�� �7�n����U�~���@�`� G��$^-V漛�%���n��1l�.���խ�Eۙ�r[��4���-�x<q�`�	��Cn����v �ٵN�n���S�g�X�G:���KY�Y�-E=c�S��@RT�w�t����&i��ݤ{^���oD���s�+3��႙O�'y/��B��Q![��e\o���L���+�(ߢ��N1O����P[I���� ��:�~��?>���q{K
�; z���[���emp�΅��c�i�i;�wW�K��;䇋(�o&�9��J1���ݝ���)�m*����@��[ÌY/�����q�G7?ٵ��ym����^��򩠁;�<�T"�8�ܢ� ��W���EKF��W�wkw.h��{�G�p���]�Ab�v=Lh�!ڹ!l$\w�wh]�����?"��Ǡ�ė�K�\Q�"�B�%�"�6ݓ�k�o���;�P���������:�Bȟ�}���d��!��j|^s�0i)��`����VfM֍Go&d>��ʴw�Kw% ח#4[b6�a{Ty[K��0[]H�v���*xF����9p�� ��O��'���흎\n��L_w#&����ɖ�*4Ԧ�c�����!�
�o$�Ժ0�vCB�U%"��Oc�F�Ha�:��$��D��^�Ҡ�S:J	��0�ЪWe��p=]�>{�iY_��`�؁;	��w%���F��0�~1	��#?��I8�v@��i��[B D��q�)������m�r#�mʠ��4��Q�Ʋ�(`lҏ|$,WrY&d�dNX��i���h�D�����V4�M �4:�<`Ǥ��$gO"Ԫ�$sg�u{M�dp�S�b-)=�����(�Bu�����W�+ �����U5��%F-���l�%�����AՎ�g5o�^:V�$j�v��g��\"�$��z���[Fߒs��<�ҕ�"'��Nak預l����� �vd�
橐Nf���	Jud"K=[\y�"�(eƊ����[;P���-�������� �Q���9vP�G֤
/����Q��`�t6
�{�#e��9E_^�B�r$9��7R���>mE�D�r��LH��Q�
9��9N?۰0u��È�-�	w˞�".U�`&����Hu}�0ɵ�ٌ5E��s�<�0%��JcD�u)"�/�0'�0����=Ʈ�d����ݛ���2��q�K0gm���I8{Q#�գ���lufU_��8����y���rs"��|y惧:
�79����ze&$�E8'����&��a����]��Q��s�Y��lU,�-~��.J֘�B��<��Ex�/��k��
fY�JĜ�f=�wn-�6\�_�T����l�@���
U�P�&�'h:���ͼ�$z�h����R�%*,�K:��	��z�쯁��	ӛ��I����)^����i�{ԕ��eze%`x� ǽ���أZ�;��os����-u M".�ynϫ4f��d��]�Vsdq�-t��ѳ����V'@+�ߚB��C�)Ҵ�7b�4��#x�I��205-(l]ˁ�7�J�y�C����aPDo�s p�)-o�O�77��ET���Yc^�}�o֧u�lP�]c[���Ɣ�4���|�H���M�o��E��#n"���O��W �C���'��	\*"`�,�ݦ�/w����E �&�3�@�"A�X���e���cMV��)�r�6�D��.��f��yQ�2����q�uYMO��`�	��B��w���Q���#�p�q�%A.�K`y���Ѷa_�<;��f$�s�И��z�~��{�u���᯲9̲]��^!��u1��|�����^�i����=��O��t��o0�3Gl�x���9���'��;8=dd��Xa�n�T��oyP;�x��s�!wPd+~[�,;kB���5a��3b(�RM�m6��a��h��B#�g�0�aPA��6�=��1��َ�2��9�8tg���6�W�=Z��bU��m8���ZH7�$�f�6הH���6���v�ܧ7P�']X\:g�=�o�}LXcM����ڝo��^�@�j�3ݵ��|��f��w������FW�r_F*	��1g~j�KG~�x�?3D�\>Û���V�[�G�KO
�ޢ}�Ń���.p&��_=.�L�Ѩѷ+�;X�����3;�r���b�=`ڃ�槂X��5�$^KV`�N��ג�bs,,+�F�NB>k�HАقY҈�^J��Ht9�����\�=���s���+��,񙇋3b�@]ܛ�C��Hc7A�����)�z�ezw6|9�&�ی �	Gb�P�k68�5�w\ũ~ͤ<�o��V�NlW�Cw���fH�*0T�&�hun��1�����;���gz[Z�[T��˲����n��+�����3i_�|��e��Wf�6�{�qf4V/�t2��  |H0�r�}(��|ms*}�qWգ��p�
æ�X���&*�[q4d�
�rim�;ō�n�rG��p�jV�OZ�dTE��)��������cZ?��п���a�2>!�I��E1Q����P��
���0�������KsP��L�����'��@�tLڧUR;Q�x�$�2���b׽V�[�L��҆���d|s��2SD�)��j�}N\�|�phwVǷ�K9��n������x�CP���y���8� '��X�b�EX���>38�q'�H�ڰ+Dxo����1yʊK]n|4�b��A�ƼO%=3�54{$�י(�HfE�S!ܱH�.M���}ݦ�} ��rS�gRXm����jM{����x 9=��� ���|ӱ�[>h���Z���v�Ó�2&�v�ZeUX��im:�1��4�]���W�t����;/`��%�RCo�)��|�[��G��YX4>`��o��?4}����9�78�8Q��:[�SY���[	-6['����YY�p�.���]3j�m����<J�]h>j}�����T�=���$�l �XZ�E�l�it'
���"9S��(����^��1
�3����9�J7E�,�������5�2�3#/	~?������d�XFC�f˞=���SJ��K� ^��=Gy#��
��7�
?����d*<<�Qs��W��~����I)'�i�E�\e}�*����]0��V�b�j�2xt�&�J��U�yT�;!�;�T�;�Ϊ*�F�ϖֺ�-��g���p_��|ו��W�"�'�6�L���;5uP�"`�W���,�
�l���+縵lD�������ٔ�\ma&�013�Sɛ�SK�\�� z�N��+4���0����1�-�B�?��
`��#�1�u�[*4��VH//�fP���%(�k�ފ�k
L�����\�c�I�r�
�n8��+�_c�ڟ-%b�|;>L��.� �d�!�z�F�%�)��&7e��Ym�@��ܖ����)�@2��;��)P�.�K7�-r�W�;,W����~X���ս#2��u1I��Yq���J;X���f>@;����,��{�㔠�'IŶ�&Ky���>e��x����"ik��f��q�9c�9ڗ�S��2� ��J��퉪6�ǿiDe9+�pۈ�l����t��-q�W���՜��ւGf�֏�<��U�2z��c3��_ze@J�|i"=e�C_�o�䗳�8>M��ڡ6�Y�^b:Q�熎ʽPf5���yӕ�8N��i�^fsm��J?l�q�ʡ՞��b�	���={Y)�����V�R?f'p`z͏�l!�^��^
a��;삎�����85�9Is,���W�5���u����l���}AB�[�R2��µ�ߠ��ې��֦d�����/)����N����Yw�@](�u�%��!��{i�F�vӨ��a���V`۽���a��-$�����)����
��kBL {���\b?S���-q��	A1Y�XG�l���,�ϊ�����LDݕ�NaFy���qd�|�=FDЛ(�]b�#�U]PY^?l��gPVu�Mo=��Q%�<��F�7�����!He@���F���y�Ť�_d{����!��`�N\K��a��<J���>�7��E�4`�G����/�~���B��L/�U����/o���`�0�<J��)��r�o8���<+�e� �O`�1MY@�2��Vb�n��MG�ÛI)����	A<r�u��^t�^�d�N<O3q�["l���,?�J�����b�ż�8�����B�tV-��T�u�V�4�(��
PDG�d�)�6���B�Cz�m}���L�yY6u�� �Q�nl����G�g)tˋ���dT��%Np���^�+V.��((��ԥ|[ȼ��=�%C�YK���͸��>��\��8��2}��̻�gyR3߬���T��]d|�����F�/�����0j�45[1pǼ!&#Ǘrb&�o�!�5_�3.��cC(v�!�2^��ET�d���������ϫ�ka������zd�4�' ,Xa�i�� BV��UY��VXQG�J� �_�-���h����ނ!�.����j�9mh���#Ǭ�)��ۂo�A��8DZ�u�'����\��͑:Є��s4L��b�U�?f���9ScZL�3:�8��G/=�-�o�fɣ��G���2��ڵ�wd�N�H)�HdAKڞQ/�TH��n�J	��F{{��(��F5Bu��y�!'�&�Pa ��d+��.�<Ѿ͋l1�� 0�����#��O��o���E��:"	CFӭ��!G)Q4Ǽ��r`���z��>s�*���MK�Ymx��!�@���_�x�k�Z�����H)?|f�
)ia���ӻ(W��d!�-�	����-��;��c%Oqd��)�w�	!���K�-���-��H<K�B�v2��,�\y���e~h��=��,o*#��|����i R�V�JH9���= 7��F�#��'	�i���<�S�ߎ��19R�Y������w��L�6x!k��xV�n�g�J������cRŌ����:ٵ�{�R�e�.���X�bEN|�ԓx�ylOM-f¥go�&>|����=ν\Sv�og<Ff@Ͳ�Bm.�+��/�"-'��h2_�i\>�(��μ���o��ƴ��pO*�{<d���I��F7u����c�ߜ�T2FN��7�R��sgr!�w��2)��:^9��@"�i���������E���O$�Eb!Кp+Gҫ�=�z��&�`QJe�ǅ�����#D������!��5���WA!�i�_ӏ
� V�%�6���k`:�c{7�ݻ��:�mg�W����VZ�De!C�Dd�d�"W�H���.��<oKP��} �q�cDs����܊b'��d��8eA����m��Q��^���<�iZrx5u���~����܎�.Cf
��R��iZ�Oy��g�z��$K��F;�k����<O�$P/ձef��K����\Հ���jb�.���1�0}��s�3��?@j!t@�C0�OK�{J/A��V�ę�z���X�*��w?W�������aj�pe9��l�gz�,T�����4��k�u�;0�0���b�]�qi]��oyEO�sU'X�l��Y]�����Rk%���Wi�?�-@4�y�н�X���k=âe����\�N{��+���B3�f����7ٜ�Պ[�6�#���Ղ�$��!�F^"�jN.���-����V�%��C�g������=n�L)��e��0��&����d�b����Ivz��<�^W2%�+=o� ��O
8�;��]ɖ�g�NX
!Pt�B���ޭ�f�v$"�� EV��r�FV����M%��/�8������!����?���m���*����(�Y�S�E���Z�n�B�����Y���bW/��$ٲl^���Z�?Q��}�)�L�����C���j&��U�a'�6V��F�R�E���M}�,�$�������Xx�����7.1݃2�Y��+�G���+>�$T����`���
�[�@/��y�7��nH�`��G3~C�D#�Lsa�Y�QC0����[B4/(D���'�#T�J8!�8��^6E���'~��6|bGz��@Y���u��̎N��ǧ,K�0.�Q�A�Oy����6�5I�S�Kw ���R�h���%3��~_���g���%�e����D_�봉TE�V�v6x)��T�x�z���"�Ǥd�Ɠ��������N5dz(`{E�N�μ]�>�
���l�E �#�b�~�u��kv�]'��C����n�k��� '��ە��*���1)=��>��=���~ea+X��ae��	�?��3�)$�gL�,8`[f��[��ᐒ��j����5Ip��1gp\���m)�b	0}La5k�}���"�$����6�&R֋Q>{D�[ʩ�+���'�gɜX��eij���*L`�����O��	2>���D|T����R3HJ����;ñ�1K���]+�y��u�ߒU�Ԧ�&*��@W?@'f?#K����V�" +�B��n��^?bRh�tMl<#u#U�~��!zk;�/�2qf���1ݺ����y٧�~���*�;�o���%O`W��l4{�g90����&JP�u60(���B?\�	���#$O�K-/��P��� )���g<�<�=�4��P�*�<���E�{�(oZ�j2����TL�{Q��`�x�c�#?��e�ێx~&.L��F��Gq������j�������d��lX~��v��G ����{�l�{Y���"Ha���S��J�)���I��ݞn��6�s۠�4[#^m*Ҟ���*R>��1w(��!�r�'؋�8�9�gA�̈́jU���_��A�t�����4u%�Y_ޥ�,ke\X�K��T��[,:z�Г�+)�R��jΠ ��g릷T��d6�^~�(���f'a�-U��E��[�����q���^��o=w��.��nG��D�S��� �V�d���o�wp7��hftB���)�wv�^����e�������pCE�A����$����ip�ã�=�y��[�G�Cs�X\�`����P���q4�զڄ\�9�)�V	��������;�8���em�/�2�|8��_k���&%<��}�F���oY��8�U���P_V�[��K��|f��ov%���G�s�ZkH:lN*]��G�g؇�yק���T��VG��<! C|Rʩ���e^��6����s�l�������<�����l��R��<�!�����T_A�q"��Xn5q1�YJ�H��vR���ۥKZ�����]�\`��@�8�+.�WR�� ~(�v��2G�UG&ޮ���Ԋ�~w5ݗ i�U��i�ZɎ.T�o
���X�̻R!߮�+�几g~�d��)�<� aybyz����L�f6g���!���Ϙ�#��!tD�˫D����m;��g{nX��L�|Y[=�S�'oQ���ص�u~���X�^�q��n�sۨ�F�mKo���	oY_��.]��#�T5tH��æc��>7DM=��v�Ly�1V[��'Q��*��6P�񎉲�n�>X��g
Ӿ��4�p�V����e�����'�qf;�G�z�y�HE/e�������~⧓��e ��a}0���ȼXhfzDp���fn��L����r��dc��$}z��8x�vx35V��
�#�.܇%�M��-�sw`��/����}U�l�<���x���n��l��~�B��ʁ4$����p@��Ul�.�w.�8Ά"�7ô<��U ����[����$"���X�&�� <�U�3a�����f@�KN���%���z���	�PO��Jp9��p߼��4�H2�e���� �ι���c��ѳ��@�0�w�C�vf����J���ԉ��4Q�d�9��`�?�kt���H_Z|�4����r-��6��j�ح�c�K�Ԟ�š(��Z��+�5d}19n��q]�¸;��]��v\���U�+�=�ڔ����Jr�����{�����5{�77N����,Yh��m�@�Ϻ�ՒU���/W�s��x�!�ҕ
>-�	�i!n�;h%$�\�8�OW]�(u-��Y2�I�1�JϛZ�͇�b�a�V[��A7����b��� -i��iӜK��Г�6G��� 1��Km�,���_d���H �h�
4���>���ӞZ�0�,�K���p��XP�Vd9Z���rv�!?ie͢N�M,�H���ԁx�ڵ�����Y��"󑱄�O�eU�=�w���V'��
��6�=�Y	�� ǎ�q��H�"6�Ȁ�sTj�͢0�A�aV^d����mop �o��Bc	�'��}��薓�g�tL8������uK�r�7q� ����(L�zѿx�C1�(יε;��I�=:�hey����Z���MȽ.��q��"FW
��Wh̺U��P�����r���}�s0���(�um��O<��E(�hN�ʲ ��m��c0�Q��GY���B����%��9r�[��ԍȷ'���T��J@ua[ԁ�]�lݱ�2�:������Ff�A�u:��n_^���g��h�e���4C򱚣�1�"�8��0�&�$�*���q�B��.T��+����4Y�e����Sjn3���$�v`��8S��?I�+��"�>�n�w^��D�������Ik�!��0.�wgȨ����_���Bw�q�j�^��݈))'5�G~{�J`̕p�XMVN3p4�����V��ג/�~䠔+��J�@o�ʱ�c�Fq;���@v7 �+�Nv�0�D"�⎋�lU�)��rȷ �C�K�o�C3y�{�����ӽBw(�^y�&T��\Ԓ��/W��; �B��cбF=�-�����N���9�����_G��������jB���n+���N!g�i�vgx�/0�i,N��ƍ>ג���IЉ*�c�C�
P����ϛ��K�R+��05t���u�/?sƜ�DDz�@����������P,���x�}"��'=���1�ӭ�c2����Z��n�-:% �2����ϻ�[S[�3]�HG��-݇�?��!�c�eJu��Z-pW4tz����J�2@#$q)�_L%a�18�$�=Z\�*nì�#8��s]C1�̏)���
5����_����C�FK�ŝr
���t�8}��)R��i�Ϲ�2g+4uɥ�����L/{�D%A
�x��w�<��*K�=)�x��l��#Éh�E�D������DN�c����(J���B �W�/���͛��t�V��]�|Yy�m��bF���ek��\��0%��hڨC�W+RI����P���%%��:�qX,�jdV��1N�ǁ�2p���� �2Ș_E�'��U�ϙ/Ge�]�[!{�n�oY��Ǉ��քqh���!���\7�oN`yw��ܵ�rņ%K��JO3pG����3Q3��O��#�����^�i̯_��	�|� z��Ϊ�u�Sf��\~8oUGS6���_ ���e�4��G߹�/(��좤xb�/�� ʃ��I����Ȓ���I��({^fAUt�c��c��h4����W������D���K^T���\�{�d�,ݠP�S���;9��j� �i
֤�|����|j���Lm��Ҿ��ǝ��,����I�r����T��ɢ�氲f�	�p�Q��]	��m�$vUC�lۏ�����ۥ�ԗ�L����cm�yh$��¶Dy�
V"|�a��%W7��ϋ@)�<��e`B*'��C����7�����8���iC6�I/||�k�R�f����-�q���а��V���n�^�=��˃yj��r>X3]�q��e�#�ELu�| � o6-�E ҕ�H�0���c����<�O�"m~g��k�MT������:G[(7<הȦ|j�٣�n|���1͢��.3:Bs������Fĺ&�+�&��U:R�E �J��d��F%�����/�n��ޅ$�������֜^� �,8]�7����;x󷬶��ײ2ܠԂ�V�Fn^ݺ�[����w.~.�Ol��eK�5_��pD'^Z�׿1�7�?Z����'�6�_�}PQ bU���h������g�}�)���cw��9nܙ�! �C��E�ő>m�Z�=3�w��1gX�R��~�a�nO[�B��=���;i4-�V���6_�;����闼��x.���,��GLdM8py���RBa§���퉹�JT�Z�?	ow�AA�C�ۻʬ�EG����~�hX�PѲ0�C̲`j��&;޲r&{�����|P�.W��=�B���}j_1��߼4�Ѓ�p�Qij�;����&٪��/g������ۺ�<�P��h��)p��DM{x���Gx۳���w��G��5��V`����Sobv ���f��$苊�VsH������ؽ������8�7��Z��(r����^vN��	���[��o�Uz�N��Ŏ������o�MV�hg�{��'�}J�J3�MoYUy��ЦJ]���2��	!)��@�5�s$ƎJ�l"�Ǔ&( �L3��B���A����i�F*��$au��6�z����g��q�ag�W}�a�g��yתtXJg�c�bq*���ʘ$x��WR��\���& ^��}|C{���<ݜRޅV�Z줐�"�8�����w[��/ؚ6Fv��sk�k�N�cд�cA�F�-���a:Tnj-3�V��@��0j����V��-�1�,w�vP��&��H���	�(��C�L��5 b͔���H� ��̢�������E )�JL��j�C���0!k��Nч��K𿍇�q��K-�lh7�W��ƃ�i�e!$ft� Zz�oi�	@�`����W*�n��1���ZH��9�˱����O��a�^�
�y�!=<�Ebڿ^��i�&�������C-���MqV�F�qD��NE����h[
�d#�6\�:uP��8�5�!Z��ɢ:3*a�n��g��!��d#�,__�/��/�{���j��8�2�Q��QU�4��fS�]����ڧ@~
Iy�Ƹ�V�Z3̻���ު.@L2!N��yn����pDl����
�Gy����x�G�k�Ei�Iz��%}�Q�h�q���F'��1��C�W��;^��l�*,�lv��l���P����3<8L�<җ��w�Sg�JfP�E�k(R�C�49k=��t��h��F��$���Yy雑w������v�<)���\�$�*6��Ų�+�nS��5v��zbS��m*��b�h�6�n+�c�Z5�����ȫ��#P�j2�� �j��sELn}Q�.�*��%����[I��Oe*H_:�x��(�ۂ��JNڐ@t�ҍb��i|��&W�w�� �T����ũgU�j�����%���� ��wKTȻuhH�bv�����f�<�Ҍ���kg�NI�����g��2��9�L�W[j~E����>�n	T+�̛�ٽ����y����K)?q�����z�g*>7���꯼IBt�c#��#<[Kz�|����f����B]��Z��&���9~ �����5Ur�@��l���;���Ő"�n k>`�}j,�L�����Nn���a���&����/���F���X�E�<4?�� f͘��%�
m̑�h�c�8�ŧٵ���#�Y��S���:�v\�L��%-s���yZ@u0|^��US
yTv�H�(�xm�t	�HҨ�Ht��P�nEN����0�Ac�n�l�<�SWg�Zɳ�s�Wp�͓��GS�5�<�d���նCfμ�xc�|e` �_3)��o�t��
1� �����S���)%|MF͇t��D��n�K���q���~�.f�{�:�1���APŽ�a��\<�P�R������u��e��G)��W�I���)�7���)(x.�W��v e$c����̲�Ռ��������_ՓM�8v�hbm
^$�$����ۀ�sw��M�>��B�5,��ayO����_g`}�|�-���V:h
�����{��NTQ��=
~�	=j�g_����W�0�ؽ�ĳO�qh�W�M���3hautG��{O�n���e���Sf�\�*?�ڦNd�r�h�����T�EGI�V�B ���֓�ܟ�.Ƥ��>���|������͘O�L"��ni����hz�	�g'϶p���˘UK��D����&U�1+��H�g�$S�ꐦ��T�K��IN���-`��T��4t�v��Z(>�o1^���V��G][^��x�����r����!�48�d�l�U����؈���?b;���� ǅ��. ��7�T��]�7��5�����:Z������6�Q�/:���N�@a+���΄��"D�S�5�%4�[N�0���1٤[M��ؕ��[�Eʎ?݋��˭1����Ħ	�~�(4�w�r���&!��01�+%��!�����*�<��uAD�\S�#�@�_t:���7[d��y��W�w!}�gi.���Ji���4<��U���*�I"��w�U��i���hٖ�2���>*v
ڸ)�)܅r؟�$�O@��0�z�9�=S�.���/Iw6���1�p)Ev.� A^	� �`0�(`[,�n	=u���Z����3`w�;v��NMw��N�&���b�9i
������-\�Cy���Z73�� ���l߸�N��[��Z���i5�Ju5@l�J�Q���60�_�e�1=Wz%��S�e�hm��;�qh8�(��Te3���&��t���w�C^�J1����w��ؖG������%����pi<�1�	�8U�I�k:��2�`���i����b�`+���RY�[������g��*1
��?��h���c#��?��(���!U������	n�"��ϗ�X�����Db�ee	]s���$���Qё؎#��w'"5����n�iW�>���0z�r�p}!��TmxTJ �c��Ĕ�3c�T�H7�]�ͣ�� �r���I��Dp���X��j*�<��'�ircE�x���Jx��*�`r2���PqR�8�؄Ő���aM=�?����H������%%A����'�Q=�6���L��D�!����C?���~)�J�uI�В�����[&*�d�_p���w~g�t_N`r������fG���V�>�����s2 s�)3��F���w"w���XG�DPF���^T���IC�_F_�P"��_H��)�I����a�,'f�N��t�ê�tnO0����'7S�K�N�(n��l���i]L�F��U�Fܭ�W21�L�Y�8�2����]0k3�|_�+Ւ���3�KE�W <D4<�B��'Hk�����+�,��l¿K�i{$r�7+�gn���c+c��������<�@��o���_&��7���W�C 8�/ʰ��g�"��B�Zڡ�ۣ���+�$���k�i>	��֢y�{�R���d$��s	� 0>S�0��%b.H��W'� ���<b���P;�7�B���>�vZ'f�l�yթ �Q�\�[�E8�cE[Ky��_��� T����e8��)#�)_�|�<	Tj���C������a`h���=r�����9�Y���� �J�;%nƥ	`�Sw�>XxŒ�[�V��3#V~�dKC���d�k�����~��z8��O�x����ޖ��i�m�b�:\��2g�̸��.�IRV��T�N�B5_�>k��h�JMK=��;pH�o;�'}N2jF�AKa�Q�s1j��"|���WkSu��쑶�J>���� 7���$"�$;��� 9K=����q��2h����r騤=Dg�CUM�WDJ����F��A�u#+��%=pAE3Ú����ߟ`��6�H<��*=j���KTNAi �9~����7u#�y��m�� �of
�����@��L���۾l�:�1��#Gy�fy��q)�V�;<�����~d��bX�Nz�yάx�����Ejt��HJn�rsMpS�@�����\�Pt�{O����ǲ��˱߯u���+�I��"a&�Tx_��/��G��W��*b�C�'��ه�n=������TǬ�W�su���U-�bu�m�.��C���w��h-!羃�^�O�Qk0�0lQ4�Dh�z6l�Nb��/�g���TZ�S��D��Pg$�{���(B�:ڗʃ�1��ɹ��g�z���f�Ȫ~�w�
U1qP޵�c4���t�g �W6�Zw��Z?`uuUD_��GQ�o�{���Y�tD�%$���S�z/�0��uXN���D_k�M�;���V-i`��M�v�	�
&O�R��	�cv,H}o]�餙j�w��-��>�g���}
F�uA��Y�ٟ'l�(|L?�˰���
99�TDӠ�
��,�\�U��1K�����n�Ƈ�gw��U_e�u'D|�8�}�#zO�r�eۣ���QԐ5ڵ��L�@<���pڜ���t��QMt#*���m\覎���UM������=]�"'y8A�p�_M*���JC������π.�齁�1���6�"�rU���ȋXR�챩c��`�i�S�毙���z6�q��5�5 �9��6�KtXq� �I7���٢��"vC��u����;�RI�Ob%ځY+���\}6�x�W{}=/�b�.g����G�ڧ��ow�+�oYq����2��)[�=[���8*t'��|`�"{�mo�I���j�����t��<Ӌ�Z�[ȕ�T�%�NƕqZ@E�Y�����P���OK�K7̀�XDΥ<P{�n�������Tsb�	񍋪X`�:�j�tU���R�d�B�'�j��'G�T8�O@���O�C�b�ʅ$�F1eN��� P�֫����ߔ}ݎ�t�zr��*-�C �����b��t<\ێ�����V%*�=��� �&r���.3��b�s�x,g���e�t0D��V��]���Pc&��b�u�v�k�,�t���䫙��Km>�\Ux��rrN���vTt�+\pW�']
� ~~��d��F�\�Ն�l0P��cO2'$�~a���g�ܛ��}���)J��b�[���?})�ے���(CL����;�բ��F���4>{@/u����?�p�0]c&$�v9��2����d���s�}y���Z}0�TK�%�  �l�*�ҼY/,��"z&\L���k=����1`#�[r��{���3�N�Y��FB�`%$t��T�(�c˩̀�-������4Aө�Y(�M��=���
�+.6pO
��c. x�X*��qV�[7�x��#4���"�.?^�X���}b�z�-�)�L�p;�vv!����_�z��UHS��V��<�zr��� �w(����4���ɜ2���Z�锥��r6a+Ōg}ZIǍs���d�b�+OB�G|뜩��|#�z���؍��i?.R�.�aZhϭo�]���ֳ2����D�e��V�+��A~�B'#d�52_�u��*�k�O�B N
�;sߢw]��V+r�)rUt�2��v/�����ׂ#_J"+or���J=���s�h��笐��gA '`	yq]���q�?��Oܳ%ۯY�	�;�4��g���� sR��jH����Bh��^��9c�p#��&՘�	lG	X�Q�9��F�͸��Bo�[�c�(���oe��̃�Q�D�K�� ��NWn�#�/���t���<���8B`H�~��h+^a��{t6�A<Fy��=���:h�鈕@�U�#��l��G����8}��Z�i_��<��߾�;����ǩmhw�K>]Mٞ��3��5b���׸&�'6�0�/V��?�͟X �ͼʒy��?ɋyǝ�bi��w�7[�ńF��o�ZT)B�u;~� F�>����s��s�FT���A�D��+����&�o��^X�p:�p�!V��XC�>t(߆y��Oj}*5�L^q�%T<=7Z�	c/�kT<D���wZ�8�$B��.�����"8H� �u�g��٨xW��_a
���b��EK�ϕ�����4G���ڈ�S�%\�1a�.J�U��Rj�\lv��fU8��P',�`rbd���v�{<�?)Z̖�_9a�f�*��<_�-N�<jܖ( ��9Smg�(5w�;kyX�u�N��R[Vj��������D�˧�M	�ރ�����I��౷����������r�b��e�R�k���}Fl��t��h�O|Z��?� �y�e�(�k��p�Ǧ ~�a�+�#R���=!��� ���+�_C�H 5�,�n�UN}�'ӵ���3��"��)���S	w/�����͚ZQ��;$�`����0��������A�u���`0�_Pu�`���~��Tn��YbO�~�߆Wգq�k���8D2����rT��k ��tf�o�U5���ɩ$^�l��!Lf�S��<�>�GjI����Xn�y�%H�r�Qe���:3�x�)��U��+Һ �>�c���e��m�<��a��=Wx���0���YYl�0����2-]/]��4%��X�s��l���������*+�(�'7�E�:��(T�7o����7� _!铭�@��L���V^#}��M��c�����Ņ�&BX�S�It��EL&�{�r���X��s<<_Й����y�Z�,���B`��)�� r�/@[�|}؝��y&��)��̇I�]w���k{�6�zҬ���XO����M�IQ�����b �F�B�j���CU��[�����y�M5f2�'�N�_U|)�^V�������|���8U";C�fb�j�ϗ�>7�R=~�L�@�4����L0y	i�����m�*ŭ�E����t��*捵���f7�;� !*�{�1����5��^.����%`��L �=����X��j'��#$k�N�X5f�����4}of��3|L���@ryu����Z`�F�TS��]ٞu��M���`=�,6�o��6.Ȣ�nZ���/$f���W�;�ۢ��^�L��B$��@���[5�U�TP�̠D�ޒ5�R��WN!�x�o:�T�6!Cݯo�����g{5�?��Q�=�v��'����e<C���A0�,��%�+���n���j�m�~��HyU���6P��A8:�EZ�>lU_� ��M*��4'NX���O\ᤨ{���-:w_k9���dR�Z埃3}�{�e����TeK��V?f��L��a:uE�mh��e[aiYi�jJ�}$'h-0ٸ��;�OB/p=���]-�aK+�߅9	�8�{� 5cx�Eؙ��ͪ�v,e�l-A�>M�6tE�^��Ҵ�89]��Հ��>�]kr���L�{�It�f���_zVK��g�!R�~e/;��Qy��p%�ΐ×`̌4���g ��!�C;���w�>��u���sk~3(�j���J��o��qI���e~tq��oZ*fT���%�D���lCh`k�UYpd�v����9|��kޮ@��rQ���̓F��p�Sܱ��.�TX0���4*�=�w8R�����X�O�?���y�*��ӥ;�������Z��ad<��'L�7�2���7ؚ�1����.���0�Q�����w'q���dr��* KZ4����d��G����3 �'۟��z�n֣y�^&q�6p`����^<^��Q�<.�I C��g�ڄ����l�	9<��Z|�X1�=�c��Wn`������8)#�o��!$��3?B�NX7Iߕ{��j���Z���βN��7�^|9�����R�{@��C����2��fTnG���C����� L�-
��Vpw��E�d�L~�����Lј�|2҉�LR���������:0,�W�m�~�{�9U>*n)�܏f�
=��3��^l����j�X�������5���6�=�ҽ���z]��L�%�%�!ivW���`ؤ�_�rxO�O�wy�-�J�&J��?g�-E��~�s����6��9��i���i������W�%��"JMO��.�TbB�#o��8�Mr	��"��"d	&�&8J'�H4j��{���J�?r�q�n�0���L�V�{g25�Tg�pI����Ƕ��^��ws� ��|i����US�ʎa�_��ϗ��1��3�2^�pi���=�1k2�E�	�=Nߌ�㞍<��_��ҽ����c����I�E���bb��M�|�d~��d���`�`1M= �Y:�P:�cpW i�ϥ��D�o���l/�l�a�����Z�V�Iam���)��V�@�қI�8��KBˇ���:2��z�nEVd]�R���
�]���h�5�������D���T��$�6w=W��x�yt��F�G�Z����+P���hA4�us�
�_�6���ڎ
fi���[��mN���b�<�j��B��
�Wir#��25����U���G0�{8MO��)4��0F|w���O��_t1p���:�(#,��O{�!剔�|����(	1ED���)%���=d_������ @?�\��Mq�6��<>�#��/ܖ�7TXG�����Wl�s	��'���_���%��@9T��
��nhR������Q���Fjs��H�`�����#�T�����k6�Y �HoL��U��_���Z?V�_1@ ��ǿ����d &���X�a���O)��<B�z�.US�=��ǡ+�w㲳p>�B���YM��������zV#0�OUǘ��ѣ��Q��I��Ԧ�<S�m:�x�
�[�P�z(��M���^��;��ֽð*./��$-���^n�]�,��2LW���s�.Xbk�W��T�6�V>w�∭ZM {��ⶃ&�n�����]�.Q���2��P���(��c�ev�9���k��`�@���Y����yI\+����川�n��r�X��#�ěc*��.�������4�QR��{���]�/��t��Z�����Qq<����0�5wU[R���2]�jFNG�Ьx��2^�����ɚ͉.G����,��K�oF��_�ްRV(��P
[ca�%s��9�|A�Me�9�L>�I=+�8�|���|��_M�w���9�o�+�g��upƈ:�"K��g�nuw`%���.��P��]�~�
��M���c��g)��S�-�h�2�O��s9��B�z��X�A�Қ����&�:�/u}�^����*��g��g@1�m@�O�+���PC��F�8ꈗ�0�O80�:��nkh0��r ���"�F���0ś�V�#��X�l;V����y��kX��	u�3�ˆvP���h+
���4�\���@�h����]�ͬWakˑxqX�����h~���4�k$��|��yᔗ�v�5-�b�ҏa�H�bU�EN�^�Ω[SR���'�|����%���M(<�4ɾ��^F��8W0�;/�qH�m
��p�S� ��O�+Y�Ռ�����&�0y��t1�y��pW�{��Y�n/�a�=kJ/Z7�o��+{7b��k��_ߪ�C
�տn89�h�'�V.���'�w� ��Y���+mH�Z>�Din�a	�1�p�?XR��f��#����=h���!�<:�a�hl���� Q:�p�i�%A��4�r�7jX�:�-���C����cS#�B��kK���^�}l�#O,j��i<��f�X��/Ej-��NQ��P[�/��}��m㰣$~�y1�Ʋvr����6N�>օ����}\�X�\},�!��ۚ�����n+�1;2/-K��2A �:E��\�-�LQ�#Wl'^�y0�G��6�2�F�f�v�$T���V�c��)�)aQ�!��Z������.
a������Zy��롷�|��%>MJ ��E��3f�Q��^��>�&�"��vڸP��P�g��ϣB��lD�	�$Y��I��[^�Y:��Z���;������W��Y����L5��M/����Y�8����%3�sx�Y�6.����;�����d�Cw��N���;��]��G-�b&L{�/�;��qkxA���]�=%Np=�������f�vmh4��A~�p��}�p��mﺑëmR���EhT��fx���p�?z��c�+9������f��=��C�x�ǔ@�Ĺ$��$��7�i:s.�_��r"�C���R_}�{wPE��ųEL��h1`k�І�w+%�@j�j��F��	��v�Nj�g�̒��O'�d�`����jM3F�F �����e�A�z*�6� ���$h��3ٟ��ZN3�ԛ,g�Ip���I˧B����U��fP� Q���qBJV*���}O;�]`���\��m�����/)�9�DVm���o��7>J�����r"ޗ:�;a���vI<����ߑ�l>���Zg)�tAG�!�kZ����m���_N�"/Y��Ђ�Mc�[���o��'��m�Z0q��S��C�x��'h�����	S8�֜����`Ur�$�w	E����y/���M��K�L�2���=j��
pTߘ���H�{Z�;g3��տ�-z��Y���21���
vg��9*G`n�0�A:4àN&B%�!9�㈨�݂��MSfR"���4�h4��A31�L�;��	�ozנ"xy*^Ż�.�m�� �wΪ	���4ͺS�F*l�����q�����Ip�bBGHm�L�iZ$DX�ul{`콲2�w���⳾*µ���|Ȩk�r�J��,��.�gdS-�q��;��������k1�[r�u�/�\�՝ZB6�p�ude�fJމo�a��,'T�ݵ�qZ�J!L�
�$ǧ�:�Bb�!>�\���5������]s���>\�I�����b�$/��jL�z�淠�����e,���.�ڒ6iT^U�!G훴eJă�K�W�O��g����|� �ձutӡX7 �ۗ�7L�|H˰�fg����)Kז�<X��ͭ��z<\!��h��U\��JT�*Y��g-��������瑏�F;c+��DR#�H#�-�Vu��#|��\1���,4s��(D�����d�.?N���m�;�+�o���$F2�i���"�G���7�M'c�Q�g� �Ŀ̓���m��Lq�>\:�ҏR�j��406�iy����4�3��[�)��.{�L���F�L�#�!��Y�VCo2T�m0x�t��/MD�-��!H��-�.��,�d2�i�̢h[� >Μ�V���H���ܡ��XwX���F@#`��ʂ�q�P.��>:����%	�g:��bRVk��ܚ|#�P��-`��m���d�����c��k�&]�G7����Q��N��G��M��[g�  =�'�MG�F$�v�&�j;Nm��E�2x���L��?۸�q���~�G;L�!$���#�����~р�-x!�r_i�b'��9f0X8e���?�Z1�)
��Ȅ�nX���0������\F :�#������}��¦h��9��$*�b���B���F(��=*��+x��0i���ƿB��o�C��*.a�ox��A_���3c2\9W��<�����r�����{�W���#6���%���[UM��\��I�h�/&N�hS�j��csoqh0ğ�QG_��m��h�2�c�x��0S���Vg�#+�;��ƿ���њ��W;%H�T�.�X�䊿�h�U��N�	_?"w֙�-���)����g��9*�"h����T��<xKޞ��|�݇����$���
P��J�J�$�;�1��)�͋\�O���x�}Yժ�6���^%���(�w1P(;G�C�e��?� �1.Z�.�����@�r&x.<�� 	��. �N��n&y���3�� �M�+Ɏ��l):;wj�M��F�3����&���=��!��/|��
ڀN�W�ƥ�(��f��?�����]�GY1z����T�mË���.��=}	���Rx+.�[�u&T+ɜ�DP�tr7-��;��4�6 [_7����T��օ�˻cv�Z��
�@������l4�M^}6���i�����
V�����A|�
�q��V�GN3ٝ �O9l[c�x�T�zO|8$��AUB�nb�����ĺ�Cv� �F�0�(���?!1����x~���h ���a�B��4j�7K�]f��tqz��u�o�bܥ�?� �(��I�j�ږW�e��X߀_z�%q�pr^1�54��Z/KZy5OG�L���uD$A_|�k3�5�����&���;���u�����J�/��u��sP� 3x&��PL,�}L�� ��7}���M��h��aVƄ��q�����.������~T)z�Hz��4���ª1P��9u������U�1��ޓu�p�KH���k�r��vp��j
�n$��S��#,7 �"pb���y­-��y2���{sPq^Ǜ��169G4�Z���S��(z��~3�P�>�#����*^��D���.����5TQ�ph��a-3���1ղl�*�ϞF $ByM:s�QY���b��� ���uf�d=e;Mf���ؤG�8{���W���z��*����s����t��Y�d :�As2����f.����������Z�zN�f��ư>ip3L�[�o���4�ߕ
V�
�^�i�|Sx��?�ii��m؅_\Đ���- ��+��0o�=]X:�j�=�z��ڽ1�y��I2����%��G[3�
E��H큫��dnQ�r���(Q���DS�.=K�+���#����r�A��s�ox�6mKR֦��,� ˡ���B����"G�M�О�*V -Ww ?�)_\�iV�f'�8o'�5����������~f�T~�1D�QR츽}ɓĂ�(U���%�g��*���_p�i�(��_��`5�P����	o\��oz�p�l�0_��n7��rjb<�6,�P0��=[��0���k��XO���(o�,��\T�b��� W�����-�,���_/a�R-��f2��b$���n�:1�_���*�v�����o��Og���Ѷ˭C��+2ϟ�Z�S�d?2�n�i�E�Ѧ��M䣏��ku��׻���k�j/Qiɾ7�<�Go���*��)�i&���ޝ͸���X��	�`9�e�كӆ�qZ�/���UƷb�oEa��AU1������Q5>1�\e�F}���|cKQP'O��!���g���	n�>ɚ���������p��Ms=�s"r�۬��z�e�����E�ߜ��j7����i&Δ�Lw���X��r$�5�Gq���s�o��(hp�#6��}���U�U���X{0S�h��ٍ/�?"�����WQ�#=�`m�˸ xcb�4a�<�g�i��~�/��ƌ!ƞ~�ھ
w�A�ˍ�lV�6v",i�"(a ��~�UD�NfR�5*@�ޒB���c�����.����"���y���O�0����r3@�޵�*B���_@4ԍj;k��$�f���IQ�6�እ�hF�ͪ��!2{R�W޾�krbk��ܤ�mv4��r{��2�h9�0��� � Q�r�
�qjyw����������!:T�g����S�l
�� ���
���^��[y�A�*S��?�eŴ�J�\���x�=� u�����qBԋ��z��6�=m�5Wq��QE)�n�%Tڶ�y���7ԏ��ޡb�\�����Q�$��%�ib[�G�x�v��_:|��nn+K)���u���	ac�^A��*�7�#� D�O�t�+a�E�Q�5
L ��2CI �\jy�cfT*�{v��_�TP�e�"�`�uoə���&��C�f{�����(?���c�¡��ԩ�#et#�u%k�TU���ꉹUg(Q���{iu��4*u�@7��z<���#Wm���&�_�U��fҖ/[��+k���5H���`Վ��l��3'���ޟ��FT;��rS�ֻ	�p	��i�Ӕ�H�C;�d�;>��^Y�G%����{!��;rw��&�h�����*O��/~��x�����)v�p����������|6-�FOX<`�e�{}5`�5p��U��\Iuz�p�Ab%�D�^�)��{��|o� ��y�7���E)7���A��bA��������r�E�l� `�Pi
�U�n��u����֌At�c)��Y�(ͻ���.����4y�G��$UB]�s���l�y�N~ӵ�R/�Q���dyr`_����[��mNf1��A�	����vG��\�xN�63��%-i��r�;U�A�>�qR�t�B�2s_�j�7k};TX1D�d��i��_q9��页�(���E/rx��Rw2�3�~��@
%|E
'�.�Q�"G[�~��:�X ���*0���F4�Pk�sh���`"����'�,����ǈ�� ����k�%�s��q�^��r���aT	�S�8EZ����Y����q�t�.q<����<���E����wlt.�����|���V��A@���K����<;q �f���@��uܔ����ShU&�'�2?z=E��\{D��-W��ua|y��B�L ��dƃ��K��T>CŦ}����:����H��)��L,UZ�k����z���4;I�k&%���C@�~K�H�B��W?Y,[u
�����>����~/���
����,��ó�h^1a�o�ǒ�N6Ї#���[erw �_��]��E��3�����GC{���;$��2���UL��jg�]"�Ƚ�9�/�V��6T�Ƶ�J����<�&:F��ȶ;��ŝk��T?����)N��D��
s^S��|��v�~A��90��tO�X���trq5Mi�+�o�#�&�ngm�>�#me�~-�S���t#�E�` �G������a�y�c(�j%�J�;���������4<,��0���
@�]��>��1RH��O�ZBvD^Xh��h�����$� �٠% �K�1"߰S0+��`/r�e���F��������Y�i���B�����J/�������Ǿ^�q�_ܐ�����N��9u�|��:�\%����.G�۹�r�L�2�|���o�B��?�GB=�d�WDZU),bq�uxF����-�&?�K��t���B�F���."�!�N�u���]�g����>Y��HV�)ã3��:>�������~��P�ZG�Nإk��lG���a�wWQ�[�C������upҰջr���������{���Q�8��@��}g#�\�@3C<��h�o�Vζ�mch�W�r���B��u듯�aL-eƙ�m�v���>$+I+�A,C��|�KX{��8��Z'xAUN$-�aR"��Y�缀oY�✩�0 ��~�Us���I��3W��/k̾ߧΐ����*:���d�;i2Uum�js�S�6�����|�b|���)�#L�@C�Ŏp�(=�G3Qqܬsy�����U����f��ͥYD���"�=�Q�Vo=
�:O�}C��$�qk����c�p��q!Ý��"	�~Ҋ��EB,]��X�`r�#�<��̏>�&\�������hKQ+�	����2^��i�L�����[@�u��Z���ڂ\���1�"��~b��لSڍ�H CQΝ狾:�ǥ��\��;�f(������'{ ����EE^�4�R*��Ui�ӈ��T�Q���־�?kWl���<�aq��W�6� sr��R�!r��d!����������0ԗ��(��lw6<^w��C?%��V���b��F�DW��>��.��h=��ˀ��FS�������4i�\�y�˻3(�XK��uX���v�_�g���D�����6{�ʏcE*��H���:�AT"](�2�P�߳��A����qm��Z#	"���d�<�=V�d�GU�\hC��@��o�'��
c*Y�,i�-�f͡���ҹ����/C:�������xrAY7X�	 �B�)r����y�����7c���ͳl)f�`t����s҄X�iX�!�sd-���M@r4�}�e�М�b���#�$����}��Z�BJ��tc3�r}., �A{�Ғ�!�T�Y~7w�����	�(�v���p<���I(V�Z�������1��2+�f�C�]i�@��U ��Z�K�H�I�s�������n��rc�k� ��\�yS�\�P����,6i�n��J�p������d_A�6��PA���\5Ì�
,�?=�]I
�ZI2���O��@5It���?�_(f�z�����O�����QK�Y��T�s�ki�b��ߍ6��LQ��Ad�/s](FOJ���ы���B���E�C\����i��Yb;�j���EA����S�N$�`��r�6Ŵ�P�j�dt��!�����h1��=�r/���`O�����,�K�.N1��$��PC���Gz�C"�:�n�w�Z>d�a 
���~۷O{8/��I�)� Q�i�W�)�]��%Ơ�ö�#斮*i<��=D����0��,9��QX��`V���M۾h�Ơ�FK���y�⑾�E	�����`�$��j`����fU����o�4��B��.��'�/!y�ƾA°�Ն�9nV���#��a7�h~����H����CMl����XX�1��3"l2������«9���-��^it�	?����ۛ�¡rOt|�����M���5"m�����>�VE��l�c��,ۮI�/˨e�G�u��W���a���w��oM=}T�V��G����U^����@��T� ��%*�͏����R@�����`#3k�+�$��!���p����fcKV�S��{�H��쇏�N"|f�C�9i�����F��&��z�������;,غ����VK���xH����7sO�K�[�dU]�G�Y9|A-�A[���w�Iu�<q?�a���J��HrW:o�}�z�w�y�B�R���<T�5�p�ý4E�l�*��' B(H��٨Ѡ~NpL2���i�֯`5������aUQ}nF��3i`��r��^��1ŷ%L�i��ӳ3ݖ�ڡ<.�|_JFA���"	��_RWl�:J;b�@�,���L�DB��4܀��'�IB�3�&�����F��ƒ=�R���&ᥫpS�&�XF���O|{�z>�]6�K����&�^����|G�Dٓ �BU�nw~$����c�S�;�p��o��6k�$kI��Bpg�1�W{�V����t�Ѩz�\ ]�F(hآd��wx���]�p��(�bJ���LZ��pK�u�\@1Ea�6{'0T�r�+�q�"\�U��(������
�B���U�֙�bp*�����A�d �.�#(S�h�s�v����~oMթ�t�W���Nٽ��U_D��"6���a@ ���E��;ܢ7�j�'pЊ�*��غ\)WTӪ��/�Z]�p�\��A��鞴�9�،��������-��V<IN��������c���4�9�٫��Im����%6���h����H�4��GJ�����/�x 1��n��1�K��q�vF&����>�d-�� �b��P�T�K��(�"����/;7 �xu������������֎q0c�˂@�C�!�Y��z�Wc��&ҘI�Q2.X�H�\��u�A���:��}��ȅC�9�� ܱ��
�����\ͭ\�-�����mT�M$��}h�ˆ�C�ő��*��\�m�!s���� ���y�&Ǻ�����\����6K���"~o����UXIv�Sx�+��WeU�l�U�۲�R���H��$&���g��!����9����x�4_���'+������<��6�ұ1\��O�V���E�ʄ�D~�D6��`aإ�����������h�H{����U�sG�A���'C�TGIv�����;�!�7٬��zZ��9���1�콐�(�˃���g��Q�dZF��q�}��|4�b�v�~�B�
�����k�7��*�:$��ă��;��I���Q6i����C]�҆VM���}z.}�:%��+��{���0t�4�"c�$�I-@�D��8��(VJSܔ�f�w9�A�X\����fFø�A;�I�<}�YxDܻ.Ù�'�#�tg�HZ����h�g��3h�)����/��Z�QeB��(@��o'Iț�®�i�6�@2���X�#&u�Nh�,����/&������3;�}=D������{�M�"N�p�b�Gv���EYQ�<�f�r��e�Dv�;썃K G(���`B%k�NmM��{�.m�@B$�5p�-��z���ȵC�3'��4�tA|$��
Ɓ�N�F��N0���;.��u�����0ݯZXm��� a�k����͑��U�r�ȕ���S]AWv띫b�!�t��׾E^�j{0���H84ڠ��C5�^"M�{��r��r����7�ĳ�)�M7��D4?v� �໥8�U���ec���_�W{�8�:G��(�@��p[Xȵ\ �b�'�طktS�ꉅ"y۵(������n�̃�@����ѫ�4Bt� ��
P+.-�`�����W.ye��f�C5�[��k��X��1�Y��G˓��F��$�	&l�wEp݈�0���}�x��-6�)��m�ky*�BY�$of:�w����tne��Sy���~�����'����)sk��� \��7	�3�<��q}E��Y@�+��ʴ^@����ˌm�#s5�De�3@(x�>�8��L����P���6q����5��;?#�'z/k��4 �`ĲZ�e�K9,-I3�M��F��e �ag���s���Z���)�r���yhۮm&����_f�pU�T̥&d�����Z=����O�%������	����4�)���o�r����y�8_;��
�z���4�H����FP�����K��q�n/n���4'X�N�#�7v �S�)S�0/���YΌ�ך����%~�	N��52�d����G��$Ij�g���Y"��Jͣ�ӡBP�*,���ڭF/:�\�@�Y_��@�Y�Z\��]�Ĕ�%HO�@� ZS^�����KA�L��Xf� fY�v4��J��3�'�{J�<��:�<6x ��-z/1�y�b��)�[Bԩr�����5*�֚�ƅ?�Bv ��0Hի�m�*�%�0�Zg�tc�.H�P��C��PO��� ��Rn�9�}DA&�9Ck�8!�]����o����:%,{��棂2v�s�}�fZ��:;�1��jZ���H��n8�Gu��h��=/�4:ڱ'�X�MAO�4�rO�NYE�-���=����2�d��o�8�v�M����fL؀�Ţ�iƟ��sY���O����3��"A"�F
'#�7��U�Cɼ��\��_W��S���)w��6���kk$hm���e��
!�Yĺi=x��"�JX e��)�#hʪ�r����z9��[M��rnŞ?��^_/v>X��)���;< �}��P9�K|-�`�$�hɟ�IQD�D�]�[wi�����u�9U�34�����������M���L�{��v�R��]�9t�̿�R��ֆ��wR����ʽR�	ϓE	�c��x��~2%�_�q�Q�@H	���۶à#VioB�|�iixlGI=�A��{i������Vw�Gr�xY������C���]Q�҈t�찾MB��r�����[	��zR��M[�?=��J^��n����.�!�@���jw��+�EP|�U��l�l���W�/�8|+=2\�4�g�h��g�R)/����������P��ٷ�S�
�ȟ��#C�1&��(&.�N0�m�*�9��2)6I�R.�$��/#�����W�֧'d����~#�IӲ���LbI�̂�
ھ�a�ې�͇���$�ʥ):3�k q�� a=�s�����\����l���7��m/��Vpݯ̛'7�DWZ���8��ߢx�A�
O8x�7*E�s,�l"�R;,��1�w����8�����	�@/k�`�A�i������'��L��J�/B��c]�� ��~s���`��-���R�֭u��+\/f�vB����}��qv´-�R'�w�����>͗�vd�|�k���Yn���N�� H:�8���A U{\��6��R�_E4�ݎu�q��9a��G(���c��3��1=�X�Ye�.�Ɲ�N.�R�P!�Lit����E�'0�?[z���}�ʳ���;���+�����Z�gԐ�z�KMp��cR�����!hg6��i'p/tl��7i2�dO@�]�^!�|Ahm� �8cΛ.宸�l��QNTv�^F?�U�k:f5N���L�Z�2\%��.� Ѓ�b.�5I:̹��$���,��d��q�HX\��:�C�� ��WQ]��1z���A�{�8\ӬP^N#~pJ��w�92���p����H`�L	h�Y���,�Aq�'�n��c���'�� 2�U@����mQq��j6�ޤ�!M�v�;޴'ܔXa�@_��璄�rك���Z6���$N�inH�ϑ�����nt�wdkH�m�D��l|Ɵ_���0r���+Q��㼨A4�2�YgWQ�BT�c���f��[��\8r�����<�?�!������n��Ia@!�̂`����T��87��]W*�U��Ӵ�t�{� �rz9�ϭǻ��	�kg���z3�xf ��j9��|^��{���"J�N�i���3-5��W	ݛ��'�-S��H5댑��Q��p�ّ��JM����p�(��#n4�[�D~v��a�]��SbRhh��/¨6�Z�=�����۾~���P)��U2�唖��C�a{�]�~�[S����&�@*9!�&X�B
w���)k|=�'Q2lw/i����7h50Cᣑ���K���i�`~i�hǊd�49��QY�қ��ռ�G�����@gۿ�p��N�(�6N˫K��p�c	��l4��¬F�A�m`ȧGۜ \�O���im�{�唛�v��Rx�CQ]Ō�*���<��:|�|n�D�;|]����Z�s.����������{e<��1A�h-�A�h��83[G����K����:i$[��i���[s�f	�$��{�W+�qz���΍B|�K11q�_�H�Y�(�~wF�@a+֧�S�z�s��"��+�d�32;֙EPaJ�Gum:�m����	��̿&���,<~��h�nˏ��N1�O�b���2o'!� �E�GB(��l�č��i��zG�c_�DWV�g��|z��pApaJ�s�������0�R���1����C�� "A����*=>s7�X2�%�:߹ �eR��ۘ�S-L�.�KM��z�оA��*N��R�c޽�Pc�2d�WSk-� �
n�K�*���&y򼺻���km�ڤI�(��R����En��]U����|
�����o	��PoM���>�B҆�Y����	lU(*F�IDAy����{�U�ef]�1�&�~�'�8e|��DI�W�lf�<��~eI�f�a�3������Yx��{GU[�&��M�l^�I�4U�ss��Dȕ�`3�p~p)#W�Bţ�P.l��k�9��l�'�fe"��x܏�9�gEw/�ҋ�GuH�7d����my�$Ǳ��~��ixF#�er}T>�<~v�f���9��n�n���h�>\Q A����������+xӭm�&�9�~�eܹ�Uz�&x(�0_����-/�k��E��gz�2D��M,�)3KYe�'��'vX|o���g:�E�ݍb�������y����1���5%���>�X�bs�V߂s��g�v�p�ƞ֘J���V�Lr�֚��D֢�m��E|�r.q�=q�uq�4��&鎸#;(/�E9��=(�F�Z��SZ2q�J��Zm�>$��K���
{o<E[59�o|��E5O�rR�xW����xaV7�$D�- �4��':7��/��S�ٵ�o䙍W�t��w.��
��hc���c�*ߓ�c�: �LX@���JW�^���8B/�7����/a��j��pU��T$Ռ��9R����Kn��`fl�Z-�b��5?�tפ�N�!2��[�$@�����eDZ�4Y��޳�
"or^���8U���|�L��q�fO#w4�z^<H[o�y�hHV�r���7�!�C�#D%�@�ӮU���vޘ�������јC�&zDt0�z�BIO�77�ʰ�"Fm����7d@�v��7[=��J{�:`��5|=�x�`D�#�eP�5�q�=�U�|
���}�4�����X��]��~ɠ�c�A�
geV]w"�sa�'6���y9��.Z~Y`+�H�[g5�em~��6�����+�ڊ���v^�u�ψ��VF�!5������ա}�Ze��שW#ܽ�'::�p\dG�@)fil���G��*l���:�
����5$ޅWq���ʫ�L�%��I�a��F���(�vi  O�Sp�(�O:��9ٽ��9�l��䀼� f�?Nm�<cX�*��&d�[Lr>��5|�����+.�|���@̐ÕN�YE;����V5�[�T�ك!���|+�H"�֛-���]��_L�K�Ϸ{���Z�upˠ�/�#'���	���G�aL����{ʄ�����}�����[6���M	���j��!�����=!�䠩�[�#�=�d3���ԫ�C�ӷ��$7
�Ru^���y�����$�4�u3�c,�'�P�1M��oC���֣�<w�
�8�ؘ��.��b)����7.�f���x���^'+>�֩��㦶i�N���i2��Q�'?�UAF� vb���Y�+�'!����j�� "��4:����`!d�w	Is��sڂ��`	����� eB�+wu��Y�XŦ��2��2.� ��2E� �U��wc��;{P]��u���m���]{�����*�J�!�n&W�(��f#(����,�!Y0M��]�I��k]���X7��(��0��JFI��<�n�*��Q=�)��;Ӫ��LMbĝ�z�=B�����6(�7�H��6l�����R����󄲐�.�b��
������\br.	#��p�cW����7Z��O�Gë��p�[����N���~���-t3��/�	\� i�1	U�罭8M<��"h��g��9X�����L3a�cM���Z�Dǵ�����xH�t�a�����w��Fl�E�m��_�K��G=b`.`���?� ��]�Rģo�?]u�t�zs'���9n�ҿ�;�}5��$R�}�C8��1��"LO��
W�y��1�p��ֽ/.������i�	\\N�<D����w>����_%oj�{"��Uq� (����[e��O3։��`��Z��~��ʙ~��i��գ���9."B��>�g�< ��ï�m+�:>��w6N0���,x飐B�`E{�8�	w7��y8N���6A�����oOM(̉PjqD�b�VE*v�%��	)^n��~�8xC�<���?�\��|Ý�1�g�wW7[��r�!)�k���R��������{O=ޤ��d���8�������)U=Z?S�h'L����Ȇ��-8=��{��'�w�����&
�K�a�`��񡶢���w�`��,��ǥH��P�?�@�**qƊ�te���-i�G�&�m���L�9����5T(���Hx�qf�N_�����X�:���E�/YQ�([k�΄VXjM�~�ZP������;�:�E�ߑ���{+Ƿ��6AJh`@dMPsVF�(8�����#�E#����E������	��O���EuWTm/��<��֟�;t�H1-�1�0�(��8%��(���j�-i�ޔZ"јٝ�.�P* v��N�	���(6|�Ix<��]ĩ�5Ku�o/Q�w�����K?<��7�D8�y"�7�+x�!���d>��T�C51����r����V���H��f�q�i�:]�O���!�HE���tе�S��Ěȵ`�[ჾ��
��m �(� �1FR�{>(���^��FA���c����b���pC$�ֲ�Kp�p����%F����7��\�f;�K|]��b���A��D99حl�%S	���6��BҏQc�1�Ǉ�|�K��i!�+8�+��<X�j�ٱTrD�X��6G�˭-����%�1d���T����ψ��Ex�B���}�s&B���vܻ����Q�4�˴v�O�h��_g����`^ߛ�l��dBt�=f3��H�n���bf���rt��Fz����3���Ox$m	R4���� >�yS��3w]��&.�;���4Ѩ�"�7{c
���*�Ϝ����f����F~7 ��8\�w����,����ɪ�񭛣Anƿbn��8?)�h�|Ӊ�|����עT�/b%�ss2����:���c�Ň�K�Z��� ȅ-��6�bߌl�
��䊜Ģ
������fԷ�i�$m��{<�ɧ�<
g��b� �;r���P��y�,'����r�;�-yŽ��GۅSK��hu�o�9���;c�&xH�����������*�I<y�m��ZCׇi5�Mn���'�!cQ�"X
�TMH��3������C�	�"���c�v�ϝ���#�9Y���rOi�dq?�C&X��e���ʎ�:�{*�;�n�MK��n���UI�'�� ��7	>(�1�c� 殂l>����Eם���)j�r�Of�C�v�p�.�ƃ�5B0(F��ՁqfN���?�6j�M��������o�{ٍx�5BlP�ugU��0�'�9�LfX�%�� so�y[7���:G\��ב�x�x�*��(5�b ���NǙҐjׯ��ce�n�(�Ʉ�C0޲ڂ��%;�>L���|]�Q��.a~h���]�Aw��������e;�vc�_���$��Z˵t��=�@#pތd�lD��nҒ�#� �%��7it�zd���ٻ~�gOOl� ����Q^l� ���W�A�A�Jwx2���NZL��R4�E�B���g�j�~�]c�~D����eIq��Z�Q�#?A"ە���d�8��/v�v��&�0�*�7�"
���ź�n��t�(<�-�`T ͉b�H#����T.;/q��[ݎ��F\��������ge��{,�8z�8��w4S���H�J��Jh�[����w>�=���Ʌ���e��Q����ύ�0K��* �f�m�J�63��H��{�w�cZ��O�/�z�EJJ{T ����c����
�MԿIt>�-f����,�͕�׋\�[����W7���w�?�\X�
�sT���V#6El�M���d�h�U��/���gJ	���X�
�G�TM0������tÊ�����[o�sO���^��L�%곓;? ��-�� Ν�A�ES�Q���Δ�`�y�bx�3({sW���
]*��}�/Pk�Z�Y����̰����>��:���(���G}�*�v�6���u�qk��m�l��n�1-�5.zF6*�姌�\^�H�W�����[N}�>�F������cөP�?���K�Qp��6yw%�ڤ{<k�;�᳐]���XƮ��<���%@S�\k��m��mT"���a=�G��w�U#�W�4���B-���ȃiP���b��霱 ]�d����l{&�1)Wa1_H]N���>o�}�`��x>	z��A^!���+K��F��X�1*yZ}��/�S��vf!neaw��L#��B��oMQ �t~����B]=|�Y�< �B3�H��1M���&�,�gZM:���^�����:��$�$�I��]E����'.�*��%0�c]���P�.F����,�Ej�!B����L'a]��(��"�*���d�4��̼tW�e���s�6,�ì<�M��&�ĴW�P%��=<��^��n�'����I�3�@U�9H�E�rj��Q����GJ��-\�{y��<o�ӄeh�����"���u�[�t�H���+n���h�6�N%��Q}�)�rd
���ԇ���H��T�G�<��pG�Q�:���/����d\INq��!�N��M&�)̓��V����6�5PCܯ�p��#t�ヽ@I��v�
w��8��	}G�f�eBjO�����V���Y�V5d�Zƪ��\1I��nx �dW}�,H����w.*�	"��p��N_��[_ӻ�&��U*~9PM�Ҏ���0N�Ax��H��G'�d)<2��Es���_�?���ǁ��);�ތ%j�^!�s��Xy���D�b���Qa���?�}�a�����GL�@�*����)���>XDX�b���~�3�}S��2ƅS��&8ͣ>O{p�C0��9��mB�`�m9P*Ni�[���Z�/%� ���5�K�"�^�f3����e�"yX��H�	��+e���v䌫��mo��u�N�7��O��^K杅de�A8���i�1�;�Q��g�X��؂�X�4G��B�1ez��3\�y,�uFb�`��F�{Er�F��
9x��(�T�Xq;�� B�\���5ǽ�	����[��xZA⹱G(��;r�����{��iX&�%A��T�!xN��d��m��-䔸�^�$���L��Ζ�Iy�<_m�ZNt|y�V��"�g
*2y�P��Q;�6d�:��Z+2�@d�єL�/��(N~�D6W�c��C���E{vJ0�x��DA}t8oj�vu~@XD�#P��/�=wZ` ��]�z�[�"���4Q�(����$عͶFh	L�W��ī�b�)�N��\Q5J?b]��z]|C�|B�����o6Q>-~jj3d6A>�׳oy%�Z���`���Ӿ�C��ֲHn�����/����ӧl�`��p�<����`k��/� vr7����
PEwzM
*:�z⌷�	�.�-������șKE1*��d�ࠕ�ԮV��`���	��}k�Y�g�AF\y�2T�~������f��* �"Wֵh_K����6T����b��+G%O)�>�h��'n>~��]����`�9%𣲱�=`�CzNi�ei�0&�����G¥���X!<�u������$u��(�R�楙K�u�`|���JX[nk�9J�5X��`d���Ǌ�y�sj�*�m������.+-W�N�Ė�E���[ܝ�<��`���6�aƳ(�G7C g�������J�%�Tv2n�_�.���7��ĥ��S��[����(������r��<���>��\�c^85���HJ�#{*U��B��R��½���=}���3��W��E:ᜎ������5!ʪ�(J9|�>Ѵ���K'F��苸��n�n:ȕ�р<)�=)������
؀j��Ih�4}�aF4�L���`ƙF�{�-2���q>����������O��}���W�Y�N�Lm����-b�g���߉�	_ſ�aoh�,��쥤X�6�	�}����!�op
\Y}�ن�����Q9gA�3��A��f��36�/����!��*}�YF|�t-�'j��Jv�d�{,�^)r���?nÞ5��^�?��t�w0�ő�)���/c�O�.��j2^#ge������g9�8^��#Ŵ!���yy���s���N�zp'Z'~�T���)�Z�Ly�o�ر\k�j�ސ>�6~rK
��fM<����O=ƔfGǮ�d�:&t�٩j���Je��B.�>��+Z��ǧT��������R��E��]X����|
��g�%y�9<v���]3� ����H�!��N�,0�����3��S�jw�-����M�XR4L��N�Ñ��2���z��d)T4�����I�5���m�����R�	�1�v*LGƁ�*�F�#|SL>����V]2 �YXg�(9��Gi�U�̴@�C6qZR�#\&�8f`r��,�"ް{��>�u��y"l �V1!�D/X�t��"�k=�)����[�<�E���o��ɔ]F�Iy�#�Ioq�t�C���t�#L�X]�o�l�H����,F��_b
� '�f|�}]o�o(:��F�ޞ���/8��_Psg�E=�q�f�@���̄�p��Ԫ_>O0�i ��D��e]s3q���G����\8����b̚��6޼��(����DD�`f<#d�*ؼ������D�KĠ�#�z4��'��<���4V�( ��'�[��TMGVK	{\Wh#��*!�df�
��>�.bG�eA�����+�=j��<���rSH�r���e�����&������;�ri���g\%�1j(���Hw{�ΙM�GD3W�"ű���P1������Lw���mNvAȷɄA3?��G��fF&?�1�=�L��aķ�pgK�Ω���=���N�Cf�Z@deZ2��V�i���麦��	R��W�����=p�I?�J*�ڡ�f�59h�jQ%��Qar@L#2��2Rs��B� E ��e<E5֪�����ᾳ\��Wf��

��-���irA�K0I��}(� L��*�B���>Z6Il���s;?F-�k�a��Į怎�_�*�,�vOΡ�, Cv����7zs$k7n�	ʋ�t�����QU��Pss��A���>��5&I��hD�oT�j��A�a�2�lD1Μ������>�]-��<F|��jw�Ñ�\���� ��#��H
/{��/�|�gr��[� {�9�j�!��N�8�zvuy]�p�4bs5'���`��#�K7�@���	[��C4�iP FR���1K��a���bFT�����lYN��A���UHW����Xb`��☮u�=�[� w.QuP,�B�&��,�0��2-\������+ɏ��ZlGS��&}�\G{h�4Qbs8E�%�,9҂)մتr7��#�����SS`�oު���8��H��?� �5ʶ���v��.�zSB1��L̝k��F�0��c��{-���	.��+���ý	�T�ƽ.�^;5q�$"�۔��j���Z�J�.���۪�~3�e��LHE:�):���?���bˠ.���p�(̯�;Z͍�/r�4�����fMhXJ�ڃN]9U3u)h����'�hf��ؕ�v43>���vг����el�K9�E�Ŵ�{�� �#[����q5�vه�l�(�j�Du${63./�Rm&r��gzfÜ�o@�\��a��|��|�̒��kQǅ*���16�~ah�<�?a��^el���/�կ��.��$|�s(�Q�nLW︂��dM��ڗ�F��,G&�$b9`A��j R4c?�r�����K� BĿ|�"�5ov�#1���|�s��B����mC�Uj���9�<I��h�I�(�+$
��r��x�5@hH͜>��D�R ��'A�0�{Ղ4*���uP)��[�"�׷퀬C����4��&�@��+a�J�(m�+����k..��Ȧ�$݃���i�b�0�kfđv#'wD��S���������8�8N�*��r&˒(X
0UH$��죈�����!XJ|�/��@���F�mT(���:�ޔ1�����!g��Q��seN��b����B���m�k�eݷuXk�v�ImO�<���>մ���yx���+DW]	�AN�uN���h�l;s����}N��c��nv�����2U���3y`0�w�xD����N��k�&oA�	�bC7e��:�Z�zz��'7%%8蒳�0�Q�䝿�1�D1�' �k殫���F�^�����'_yl�1���aoD1;9t���C��^[ "yZ��5�R��i��KI^���I.��CU�F�B
L��t*�v��W-�9(֖0�	O3k蓯�ߋ���mm�d�*_PV�Up�;�������HJU������Ą慷N-R�	�������|�ّ
�G�v�r����(*l@A^_
L�JPn��뉩]�t�m+��
'o�������eEhalb���/(��*��0��9u���
���oM�[��tL*�x�l��`q>�Ǝ��X�w	�}�cg��Ǧ(9v��}�w���]�1b�}�<����<�Q�T4x/o���pk	�њ��q$�Wȁ=pK��}s�Q1#W�-F����f��pԸ��,lŊ�xf��&/��Gd�9��ڥ�9��H���`�}��w��Mf���b �J;)�{��C�`�rZw��v�1�_�\��z�{���Hˁ�$�,^-N�_e;B㣂X5�m�V͜~A85�;���nz�v�Y�:Jd�!2��;�<j����Gr>zW�fV��3cG���'���.`�>�	<p�:������Ӫ(\�)+���d�0|n�Q��ښg�#7:!����yV�.,�#��Z�;�MKM����i��o�T4�ss��$�ۢձ&����E�z:�M�"a�i>F��UPPii��AJ9�tvW�o`����mQP��1(�伣�'u>��vT��]u0�]\�'�^nF���0!��,&�Y���A����F5���������9�%)�����9��k�'-�|���r�l�Lc��M���1�K�
��e�D�k��&!��� �����^� ��A+"�f> �R�8Υ��e]2ޯ��V!��Kf�|��]J�?���\����m���y@���?3f#P��l�Ǽ��p��~`����ݤ��z�N�4,w���ǎν6���F�C��t��`��,��a#q�����0�=���~1�잯q����B�ؽ�|�x�O
+�/[7}�A)�֪ ?�$=�U��
��1�^��Sf�w�)% �HE������T�H�K��>��fT�aV@�8l�e��k���|xC�D(d=ࢫ%z��Ճ*)�uC�FKԻ���8����ÙB�ʩx�
d��E1��/i�ϷA�aݮ�mCUv�`x��D!��qe�}��E"��&*���+��J�s��T�4T-0��rĽ8�7a�,���H=l?���63��+3������� - �N*Uwa��@J��cz�E�,A	'�pF��m���8�tJ�-��e�i~ĝ��C�|��p�;��t��������)�&֎�H��9mx�gٯ�m�'0hN�ݕ洰yÛC`��&��Ǳ޺4��i�H���𥿦��R����� �oM�4�=�-��l�f��G�
r��4�B�;���	�"D���}Tl����%){�SG;:,���OJ<�M�-�u)1ʝ3��h��s�_��Ƣm���)jc���$k�8��s ]��P��i����,��_[�R�'��l�}���c}�m�t%g��:�ª�{���Oe�Zx�x����f��1|A�D�8O�1�ݬ@�.�v(�G��p7��p���߹zGFP����=�j3F���!hS���-*R�fw=��4�ƹ�|St�Ԋ�Yg�o h���\��e3��Z��6;��h<@c��kX6kz���R��d�Hz1�����2$��
�.׹���F�s�5��W�0v��x��*n��r�F���{n�W^t��c�l���:�+��'�'yg��X�<�s��~-�
䞢o������֨w��Gw=3�8����D��(~�Ev*�r�����>���?ˊdC%��c&���L! ��c:]��ЁaO���|��BNl��r�x'��k�р`-��aV�[�[��o�HvY!,c�@IO����eöR�6`6�*U�A��}�<sA�ռ@s��M�n�m�j4�!+tX>��2M�v����
��srPV ��v��e�[PUG��*M�ؤ��c��5��h��l`;��ƏA�����sk��E��S*�2�ǐW��'�dR���(�A�W�9*-��ɋ�GIU�r�u�Y�5�k'�������u_�B_����)�,&Yaz$O�y�E�"�F�� ���õ�z��(FP�#c'�cb�D�������]{ĩmav��)�)OY�o��R����(AyC�*�#��+��@g��3��/9�^��ް,g�U�F��<���7��:G)rq�c���*���31a��sI��j���6�)�H��!��\��q;�]'bԣ F��� }��	���!���m=�4a:*T�G�Ÿ/d/C���'رg�J���Y��*�~9f(��a�1P�jO�&�<&>��VΙ�Ǖ&�V,#:���>q�� ��{�wcs�jA��>6bǋ�7��;_扰���۲x�P�&{5��)}#���z��MI������I��MT�B/�<�ܧ,��̇��'_��Y��Nm 1�+m�"��_n(W�ױ�j���2b���DdX�I�6�q��}����,whR9�����O���'��V'���*x�Ά�o�k|pJm�����oo�o<0�I��A��^����pED���Es������<�ǫ��9�)�ߺ`wō!:r|�����`ԭkRV$����������R@���~�%5|u'�C��-��>�}�W,�G�K~����3�S5Ny��n.��vi}�q�k��=�oףǛ�X}�R���I�Şc+g��}Ul�h�z��/Lg30��y<��
�EՎF��Fc�bp�Qc�J�����Ňz�Iv\˗����/(Q�Q��{�������~�thw��C��Gwy�9F�aՐ�(�`\}
ɰ�xȵd�;���	/�$�Λ��� ,�6�&4&���RZ�U������o�*�Ϸ.Z[vN*��р8\b�~�"\�#��~�Ƃbe�g��y�)R�':��iN"��/�#8)�t;)�)���m�>����A��O����b���~��F�K\����l���~7�^nUdE��|�DDz%m0�
�u++���ѓ,�������N��1��@ŷ}��J�.�B�;����{�^
��4���xؓ�)ld6�P��^�HEP��o���^Bx�z��%S��^2���`}�����?0�s��-L���(C>�E��nݿ.k�e��ձ޿/	�̲�U� ҳ�]mPa��~�1�"��S�Q�W/����z	c*�����Ĩ������l1��F�7l'�������)���UYB�Ĥ�H��L"�u2�`��Q����/��e��8o~ܴ	&DS�+Tp�����	3��X-���% ^��;�������0�D�n�`4~s3�
QEࡱbF7L}�p�[K�W�1[�8RYq����B8�sB�	n�6A���ݷNR�oJIAW�v����?Ā�1�sE����P��$�����G;ч��PkT���.�eY��0RA*@��S�Z�26>�1JڳƎA�c���'�'��G{}�o��s0|�K����o�R�>�  ت��V�2�"��K��V�˖���c���ZD�H����ƃ�R���nؗ��j�^
T���1sqX�/�c��~x��y� P�@�de�����$�h�)A{���R�V��*R��T�����}�<�E��:�ĈwqI�jo���|S�qcb+�i1�.ŵ���u�"�"�-u�h���m�d8�O�	���i��Z�9^Ļ;����<�GΠ�p��9�D,�\3i�l������a�+Ɋ��O��gĘ�
���zB0^NH�Ϊ��t��"�ղI`��kU����ԣQF$���0���:D<r����q͛k�$�,�~�o�`�������7$.,C]u:�u�������E����( >�/���T��T�)�6�Б�%%]i��R09AT,�f�#��8�p�8aN�,�ç#��,��e��
09|�Hu���� �_�Ꟊ!,�$�m��"G�WO&,o:�ҷ"Ub[�<
Z�������~�E���H�y��ۭm��L*�/9J�zQ�H���j1�&��kOA�A-�4cE�M�d;���&�]+թˀ(�3��B�L]����C���<�a��^�)8{r&t���Z��)d^N�>rh�%�_�x_����p�J�~W#��Z�@�[՞�����7��#�9�=f8�ׯ�$��J�r��rI��$_ > L�硏���@7ݻ���N燥QN�����HOҕ�����ʋ�f�ٷֵ���F&D�M��D��1 �	A��Ĺ�B����&��h)EHwh�Z�������/����h�4-;�-�{��BA�����+���o���_�7�'f�K�����\��*�@. ��-hA�uX�M� v�30T�U�����9�Xs6�cR4�F�1��廉��Z����4+�CM<���c9���|F��8k���+��˱�=��'Hϴ�ؕ�\|����X,�uޙU�`I
h����4m�T�����&V�2�����M����N�\Q� vH�gx�e��*Ҍ�+�[x}��zXH��m�����]G�ֵ+G��=त/�M�-+�L�;ezi0v�\x���݀��sZȨ�e�+|��ҷ�ʾ��m9������D5klV�Ʒ�(&.�Y
��n�u��f=P�t��Qu	��B��:�4��+y������H�ĝGm�Y7����(����[xE=^��sF<����6v�k��7�>�v�z��J����� �[:�jAܚԅر�����+���u4�%���Um����~0WN�T5m�����6�����vҊ~tf&Bm�U/����>u˓�����cq�~��Y�f*�Σ&R�J35@�:�;qq���� c�ns�![M�wgE�ȕ��/,�t��Ƶ*(yй�#��$���v�*�C�U�IL��?<�:����֑.{��d�q���*���/�׍O�d�O妬H
��V�A��#�(#�bO��U�1��\���m��?� �ᱭ}=X֊'X��a�S��.kAS�m��#+v�|��Up�:�B�h?y�'ֶ����
��OR�׳�SK���	�b
�T��eE����i����J�Ķ�nO<P�r̳���i8��%��Iڨs�&���A�b֙yK?���:� 8/�H�V��)�'U������tF�F@7��u��u�X���e�H�D8!.^>8���'3��"��B��d�+�0E�?���_���
�(mG6����#��[��c\�R�|Kk�H��!̘>_u�r$�hIŕʄ>_�b�+ {�8�T��(��T�ȿ�e$=�:8-��U{;��*8sÂ���������L�OG��m�tFX�Li�i?�>��$ė�O-�)��T�j�������<u��������J��$�ԴcǔFͪҢY�p��Ͼ�5��G[�4- 	lS���=z��7��8@�� Y*���mÌbB�R�R~�:�������{]�?`5 R/�G�F��W7eJ��G�6���:_�󰬆h��c�1��5+��4\E3��ڐ�*e3�j~D#�ن��,���vb%{Eӣ�����N��#|�)�*��;�k��K�h�=�U���$��-�7�XQh��>���|
N���;z�D"���L,1&v��=I�R���Z���-	���g�ű�s�[�b ���X�Y�[�R'9M���`����̂����ݍ�qm�F'}B��;������S��8���m�5N	�(�� ���Z7FE�c��i��Z��@��1vb���15a��g�	�j0�W���_����*�mk�V��
0��&#���3�K(T��bS;Ū�cZBb�S:�*��m/��y�0~�-�Y���?��ɟ�q_Vm�[��P�H$W<Yo��3�T=}MZ�4K�c���i����Xރ=XhƢ�pC�����u�KC���f>�n���u;��{��ٵ��;q�m�«��1���1џ��~Rk���ٶL��cd�>���b�P��%����d�=��N|�N��n	io��m�Y�GV�tg�L.�ㆠ�Z��A��_�2���g0�;�(N�G��L�q�՛�|ta��%r��+�Iݎ'��_}�E���+�"\ �8���~�i�8~G���i�Oc}�����0�����\�;�v"�����6v��M}߲H�T�<e!#�;�ִJI�n'�Q���������ג�7	�W�L�"x��K[2�G��/���B)���B����Y�i۹��ic�/���sz�>'�L�iz�'�,l#���P�/gb�~	�I]5HA ۆ���/��c���JC&^�3�"'�� }��I�o�±!�b	��I�C��),�W��2!���x�����}v��N�?�m#�A�G�д�K��P��J�xu?X�*�nDD!tWZ¤��F��6'n˯
�i�ꉾ��kv�-��]�6\d�r����t��y�,y�lrB��s-��
�:XPS�}(��r�f��[#EI^�	�k��9Kݴ�/����0ƉݖvA/�e��ǧ������ �y����q���w�y�Ϙ�K���]���!�Y�w�@��W���A�����ӽwv�C�t@��5]*�Abm氣�ҩ�������y��E��qzw?m�qrG�B�ř�<(��ݏ�u"Dέ��c�wz;�l�X�)VNF���Uު��y��׆i)����ᰩP�?a�/��c�EbF����������ȵ��$��R+c�\�L�{�N�Ɩ*�Ȧ�A�EEO�ƚ<��q>RmJ}�m˙�b�ȁ���%�G���N�>m���#�����|���6�s�VB;��e�-_Մ����z���,�����ubaA��/����9!�f������A��O�YR�$Υ� �z�Izlz^�����ͣ[�1��L�r���4g�����I���X�ji�.ū��J?��f-�ىȎ�GJ�R�"S�삎�zk#{�!�ճ$-��Crt�]���='�G��:7"`iP�;�%�C�t�!��C�!O��,<�~�N�L�����%��}��6n�T4�x��9��[_Q���؄l��]�:A�+���YJ����6~Zb�r��`%N���v��T�"�������#�s�p��/ocFk+�v���6s4��O�d�*9�1��HPZ���b◇.�+����H�P�n6�+I_Y�c�p=ּ��[������
�gJ��������y�������Ӽ2������F�W��l�MJ"�D�^���^^� �[�K�����t�m��жg3�@�\]n��#ૄ�;���}��)�T�?tj�Qԇڏ|+�Aepw�N ��4��u�U�?�F-I��������z0�љ���d}����}�O5�e�t��vI�Z�'~�����I;�p�,��u̻�γ��.g�����^���i2�dߨ�!W�����e��H�l.X��*���It�g���W�>+���1q�ߒZlb�JG�G��Z˝L���	��q����K��R̥�6�ϒ,v�Ȇ�(���d�?�����t�(�ُ��F�]� ����]Vbp��������⾪tU�?co>n7c��5kk؎x��d�.ɻ��K��uj�ߥ�A����;�t��qziңrR��|��B�@׿�72�M',�E�99��U�y���QE����������-������<��O�)���Sʂ�CQ��8��Y�t�h��Й0�A���ǿ�z�OZ��bʆ{t�7�&��J�5_�$W��3��TV����>�t��_CHJK*�h*���U9�F��[�/k��y7o
���d���� F��q��P��X�{TFR+)IVr{�Xط�=j=�3v"1l��sK�L����T��ڹӃ���
��0`������A���Z7	�:8|^�@��oc,�����3@	H�R��'r�6���C�Xg�+�ڤha�n�0�
QH�j	��Hn�P�8����!��w��)���+��'�W@��l"y�Ѐn�B�����ņ�	~�IH2�M�G�&sd"��$p\%�Q���yk�WV���΍I��)7��ƽ�����g'�uޔX�v�C�>Xa_I�D˷A�I����}��2�-.��	�	>\�I�h[��{Vv�Zy3����4��LZ�',�܁H�a�P9�.��Է�@\'�	P1晒���>	�F�?��OC�ja�a���'����F4&~�!z��B����z���a.�5�r��R̘�<Q��\�vr��w�gf���Y;"�A��K�|s��W���s����Z��	��z����t\s��y�7�|j�d^��{j�p{��/{b+�5Pm"�߳JR3��$f֙��5���φ]NH�]7���N#2����G�%��mb��5=?��.��e(�]��E�D��)����y��ہS?C��b�N��[b�5{*P�)�]��[�,p'l�Ƈ�<�7 )�E6<ڠ+��ֹ�����5�����r���"���H�+�c �=�VU�ظ�LQ��FUb�\�n�� 䏔�W���膸�E��`�Z�b� �DS��O��C�x6|�9֘��8y�����K��!��e{P������Z�gN�Sބj��[#����~���d�v�T4�Z�T]�Ӿւl- jR���P�tO�Z���che֢���h�}��"�� ��~y[�l��#��7�Y�?����C�J�U)��9ؐ�٧O��N����lI-|�mg$*�{���8)���\_�g��Y�U��T��O�d�}U�\!j֎J!Q����mn�x5���QS�7`g�<�~��5�@1��,M�x��tj������	��/��+mȩ���S��!� 	>X*�Az%38��3�4g"����.�7��ǂKȓ�A����q�%G���M۾Q��pg�O��N��*�,�2�^u!x�ɉ��	�J���o��pR"�~��V�Ѯ�1TbK.�_Xg>���	O��g+���'I�(�}^y�x�S�����1X}t��y�S���!Q!xg7g/�ј��]����|-������tC���<D�ӷ�W���vy��x��.5d|�=�D�����v����~��o��c?\�KA��oXd��q"�\-|��1_�h���Kc�?��O��s
���:O�,Ƽ��4Y��8�!��
����_$ۄw8Df��:�3�،z�e4��i�"�3��zQ���GV���hM�r¬��0��}%�CKsAptP����}�M�> �>��r�riK�~�U�K���ˣ�S7dr�t��_�oq����+�8��r��%Ȉ��]M����\;�Jq�y�Urg(L����tM�M� �SL��XƃD�;���fe�g`��8�[}�5O�#��ڙ��3õ	ԟL�<�0k'���u5�F��Lv�%T�X=�^�_�)5$�#�ᇋ���)����+">�'�����H](U�_�&�3oGr�]5'4c��f�:�>7L�L��b(H��&J	�ID�S+W�QM��z��|�R��тX50.D�<A��"[���=�N��í��I�)���L
�묏'h�׍��
�����r˼V���1� �/��ojöo��W'k��R�&x6��U֩e>�Di��Ϗvժ֍W2��S��,+=<T�s�'��ܞ�Qŉ�o	�����8E[��㚼�~�S�����ހ����J������tz��۝.��*G,;cW�d��x��r���F�V��	E���
��E�|r�%V�I�+$��k%��~�ω���R �����{Y���b�&�;B!�1S��*� 0�NQ++ht����-s^ZT�Zx$\�@����V.
N���t������L;�H�j��5}og����(r$0���W'hd�l]7�Ar����PAEs�΄w{���ܙt1M���k�����	����jms�>���ض�F=*?�Ax�jk�l�H���up�{���nj��@j��0�)8�0����gYʧ��	"�( �8~x 
\��G�ka[Y�Jp��/S�*2�M�>v$lQrƵ�w�*��5�]jUmv�q�#5��խMv�QR�6s�^j�i�N@�7� ��������w���>�.�[�9��+i7bk����"���,���B�k�I�� %�b�m�䇽K��#��5Km��g�r�[�l�������� �jY�_�������7�����3��yH�0�%A%=�4�8T�:T]g��a�1��Y+�ך�4J�k]Ц��3�?q��lo�L�z�.:��������[\��^o\�~Y͆�����i�	���3}?�y=G�Y�-v+cd/�1THd1ƞ����s4���ڛȤr1�U�-j�$�"˶��JJ�E�ף�ï����7՚����DJ�	��D�.eR�{��ȵM'w2uLރDBH��o��h��~����1�ȵ�G�2��=�F�5�.0�}�2m��V= ��=���o��o9�Rwvܢ��)3�ap��uاNSJ��m�2�ؿ.='���w�JNA���ה ��X�����|;wp���͖6�r�D�-k��=6V6�M��������·����K�33�R��D�\7�L��6��?��U�)g�R����K��Ē��ة��6c�bM~�`G�՚E�i�~&�Љ���7�	P��u�{lM��P�ñm���zG"~�`��	O�q����XJ���Ǫ�& ���o���c�����6�܎�]�x����U�pDn��8à/'9dd�o�z!T��1_P�v��V��[��t�v��.?6b�Ef�W�<���P�R� p:ͥ=���D"RSE]�ڦ���o�sW��J�$�^*����9v��KhG|����ߑS�X}t6h=].�)6���ϸ dc�ì��3,S_�!ϯ'�=SX�)X�A�ѹl�JIW���H��-B�^���f��]�4~|��ߡ���j�H��s[Ծ�A�:d?�M��xЂ��텪��Vx�H��ͪuWO��w��>߂���C�Fr8=�q��L��oU�ٯ�̠�_�l��x��ګ��|��F>P�G>#Y�o���/q�Ȼ��Ѣk-����w��6L�e�(����!��e�z叜#\���؋:d�7��j�.��㤒�t�{��iۍ���ܫd��=]kjWd3�[���Z:Lɤ[Z�r�?-h*3���m�mg��ӕ�I������[��y�:D�q�/��E5�u8�lg'�|����%�Mh���-i����!���,V��\��k�ֵ�T4C�m5�dN����ۥخl��O����=����˃�Cb:C:��y8^;����0�����9\ ��x�|އw�[R/��̈́Pׄ����'��C���u~�`��%�g��t|e��r^MS-fԔe]�(��o.S/�gf�>���"`-���m��j�jQKߺ����f������2�������	��/�G��	 ��c.?c�G��oc���jyv;|Y!��\�"���\$��q���H�z� 5�^<\w �$3�Z����ks3ZD����ޯg� 	�o6؀l8 �z7�_�3�,ȭ�&�x|���@��y��} �Ja�����Bg�Y���S�\�@H��@��x�����Q��V��yQ;��T�05rug{v�9��A ��議h��jư�za)kM��Y��j���	�Y�^��/�N�ll���Xr�`����님������>%hۧ�5-�	�R>|D�O,p<>_-xB�VZ�?��,�֥����H&��J�k��.~5~ p�S{�O3����A@d��P�,��d�ϐ�/=��aĦ�s|��OC.��}�]��(�)��Vlg��<�P6���4o�%����q�CeC�%�@>�9��'��VH�r��v�l%b�b����h��4&��C�IS�
���1�1�Y�6юgMӠ&��Q���Q6�\�\��?�m��PGM퐉ɘe�	��1z^Ψ$-+7z�R
F �9֗V����~R�.+���^,��Y�\=qx5�����A���<T���,���xgO\f_��HGP��(bG<�	3�t���h��L���L5p��G�'�P4>�MN�DS���]��=��Q�������(wfon���+�ox7�~�U"�]���'�.G��]���l������ބq_�Ƀ�?OCQ|����N���s\�c��	�g93U����~�X7�=��R���8;\��x/P�9���D.S� �GP,�����m������E���ԼO��ZX:���%3�e�QO���˨�Yz^�����v��}����$U��3��Fǂ�&�i��a����m���Bop)��~3I�:�u�EGx*IY3�wo
d��G�f�܃���1�o�aN(a�H�2��Y�#[���F��|aS80��[7_i0h�)c��Rļr�q��p��u�)���ƱtD�d`�M~�GkƤL�,*v�[��(�#�3IN?)�k�(k��Xڄ+��W^�|oS}D��˝z*�!Ǿ���]T��2���x�W'�W��k�Y�p�%��pҾ�3tl�8�'�kzYB�oց2��'��vJl[�����p=~�!���Fd�O�)�Jz���y�:���	������3$5cC��z����9����
��=��(M�2Š��?��o-B%N�	(���9X��g=�m�f6y���9��G����ȹ�}�r�jŁ�;r���Fr�k(O��R�0�q��\�h�I���,��K�ďs�R?�4��zV����D��*���6��k%.�G�W`�zA"iqܱ���'k�k��pH�K0Im�a�(^��:ة��8�9j�ٖ��=-:��!�9�k���4W'��E�[e������V�\��[n��}����2,�V�I`�U�����#�S�݌�!ĳT�H;m���岞%���������k6��x���Va����*��z�MI�9�S,�u.tE���Z`(���h�v2��E����l�����j�� A^���qCc�s~�~��~ �"X��C;mVn���+���6����կ��q6g�h
Z�#���.��`�^���� ���vhҮL�'��RmSKm�Q���4nյ��
ˋ� #��3�9�
�5{*����h���14R�I� !w�Buh:�d�ώR��������v_��mh�w*N�?��rU�&w��R����0����l�x0���S`29f�N�uI�m�:!�e�����g�=�8Xb��J���P���(d��+H�	��0�W�!��b�=I|��ex^�W����̷����aՎ���
y[�BN�b+^5�} z��\�EƲ�_����a�~�d�~��0�'��N[�� ��!�/�xI���;?�>1�kBN{R�!�U	�  �w��{����H�� )t-lQ��W��/��˔�,�\ÍV(�Y����S��]c��.����շ���=����Z]]X�:�w�!˚{�eli1�˖c�[��E�|�f�V���X�]?kJ0+�D6}A�vN��Z�Cum�\��tY�-�p��U�S�@ ;?O��ŴdI3�2���^T�ٕ��O�Z1*��%�~s-d�+U�Y�I;�r�U�F�-�6�J�H�Pχ��vS��p�%�JÏ��K��{{4��ؖ �g���
\���F��ېx�ΐ�L�0����>����׫��p2�Ip������1鿩N�:6Mt�}<9is��`�w�Rp��nE_o	"hx�>�V)���':խ�}*m�4���x��j0)�W2!�q�]̣Ap�����JA�e�O���<��eR��s<&��
�P��s���"oI�B]d��k߷Bv~i
�I�ME( ���-�|�bT�����'���+����PS�3%��hX����#*����O��MԖ2�� �U�d^�5#��!D�1��\��K�̟�WP�H�8.�x7_\��-��%M� ���z&;����z�ؒDMPu9��p*�2����G�*��\�c���CA�7�D�dᯨ�Q�3�9XB���r�����ɠ�CW��~�-�R���:U���SYy e#�p8P=ioV�����	?��V?b�~u�<5��BOځ&\Yj��m�]�p�5C���V���e���Yi	� ���R����G?T���T��(E�]IEF�\v��OKEYl�b$/�� ��_ԬżL٢ 2)�G��GMg.����#\:��c��,~����%A;�f��@~�J��)��:Q;ҸՇ2$D/���^D����(���������$�R�0��~=��ѓF1H�:�w�2A�~��s�ri��e߹���Z��T���Rdz_f(��͏�x��|8���#Y���]����_ϯ��R�Q�h������!����u�ئ1�#á�Y:��0F�9�	~5�z�Yl�B����I�!T�K�qKJbK�$_�e炴������Y�����%��T_�1�I�Ɩ]��e	%f�ͯ�9`�]��7������me�r��$��v����4�=�/��	�%�T�իo.�|�	��Ŝ�e�]��ָ���mܾX�0}|�z��F6B]�۴�?�ݴ��Eme��(���I�u7$���z�T^!ׂ '|Z��o�O������pi}�m1�T=p0�K:�ꡬQ�PL+�)������G K���R���@�ݠ�v�xq=�i���R���|�-�澔��&���J�[A���\Q�����F��L�?�EY� %�)b&�w�Caa�<�7���uw}g+�GT�"�[v\�/���b�)И�N��{<�� ��Mb��B��`N)Ǜ�}��7�~6�f�[�50����P��_��#�R��]�SP�����g�g�;�C�[�>�!����aA`�jk������D�u���7q�����I����Vh�&�ϻ9F�k"U5���q�j��Ro43z�Y�a����w3�{,&����pJœ��ּa�y��b#�Y�-���|;Q�0�h�"˅�=��c�������p�����9V�s���Z?����X��L�*�6���%g癩�U�kե&�[�_�\_eJ��A8 �J~�F8���V�����gN�rblm�NW�Q�`���4ۙ?A�a���e���;
�~���S< ��M2����z�����rW���PO�F#��G=P�g[Vm��!��qϞg�գ*�[!U�4y��
4d��ֆ8��Z=e�u�eb�8)�kN�v����­/}23	���MS&��98O5�{����9����n��9�Q��^PMܗA��PNYq�D{�8yp��$Fqԩ��=x�%N~q�]z?�	&��+M���Vg�4(�nT�Z��hJj��ꤰh}�(()M{�,0X�0)�'I���&�l��l=;D��2h��Ǽ¾mo�c��ks���qA@Gh���c]�m��Gǘ��l�9�?ϓ�L	��7T���^��WՒ���Lo�� �}�h��-zF�U���s��(��S���? �@�&y!2^�Q=��^�d>jA��y+�Lf,y��,���O�� )�XtE����㥿�_Բ�O4J�t/��)�D;=B3`2����ޠ�%3]G�@2�^=�@&,D�B�\=�L_����O�A�"C��"ÿl�s�ȕ<����p��8�Ԁ%}�ńY@��ͪ�d�@���&)\����q�T�q���2�^�N����a�F Ȝ�G[l�;ܙ�Y"�-��u)cB�<2������u�!BY��+����bIB�oޒ�1_Ya�xO$Ԉ�)	n�_�������S^i�q(,���&t̒5bfeM�B�,���`�H��[�:�ikj�������@[A�J��zy�QvY��y�Z��� �,�2F�����\7�%uY�����"��{�W�nHƚȿp�-��GO ���".<w?!��QbkJi��s��B��_*�_WJQ(?�S�����"���m�mP���A�	۰�BC�F���G�o>��е��H�K�ɱ���߭����oY��CǸԐu��$�Հw���ʞ
h*^4�m�NWIk�m$r��:?阢��`KvsiU6Ȓ�V�LA�EO�����Y�pՀٻL)�������
� �����}(�%=��0>fc��Ȳ�'�K.�(�8��֪��������:~h�F���.)	�	i�b,Ӱ��[�]})��[����p�"�(��c�L\+��A=a%��l�K�pnX�e�o�PS�m������kMFp�D}�^��]�U�����C��2v��9)yM�S�A�񿂸a.�󴗦^O�C� ��c���` q��7u>��fCI�E{N�#j����˹��i����;��~K<@�e�_�.�%i.\i�vEy�._�d
8�LT~�,_)�$��
�jv��kP����z2l�]�Ѽx���lv����;p�,����0�M�̕�&�h�+ď���z��?]o�wy{���&,�K	�	��;3�w�;x���<pPۤF�����~x��^b`�|��������M���0�P�>�3��K������G��xC{k�6�3��9��.i�bUo-+d_�Xz�f�Y�tH;,qӼ �jS��h=������U1�HWH�8��T̟U���J3 V�Ԙ��&^����5^�$��C�����j_�PZ��ז.�U�)�6&�5k���u����IV���64̒R?����?����h�[��4���Hx9ukY��Ru��3A�6��U\-���S %�,{
N��CR�,i��ʎ�"�lbL�����n炸sz���/C�.��2��~��/na�;ꝴӻ���{�S��Q[��O�(�~������~�n�*�e�RJ�╯\ƈ pUT�5��u�[���tZ19��g���V��0�tZ�n�i8"��`Y�x3�+F�^I����U�����G}R>r��yL�g�c��d�W��2�L�3��k���+䄧	���,]���C���+_k����Rw/za��ڣ�QE@ՙ��J�Қ�?F�-�7}�l<e{�!z����W�s 0�e_�{2Ht�R�"��W&�Dq�ד�� �=Ff��/��w_C���>�i��lz����\��%g�ܢ���s�rL��lϺK��J���Z����珇3ma��Ӏ��%q����ӳ��2�a� %��T|��e��1������N��d�I\ �����&<i	�5Q�:oP�-�yr�0�4f8�W���ch4/�Q��9��&>s�s��_�=t��&�_$�k���J?�.�ӟ���|&��g���ذ<�8$Q��R%Û�yM�DM)�&;���A_����]�[eִ"�p{��R=�:���Z�U\�R��^��*�ގRP�M��e������;�����]c�َ$�5��z��Y1tL���x]�F���8����PU"�BnzOz�r��%�W�� D�	��h�t$Z8F�ܰ�����h5`W��_�������O&V��j{��m���Lj�Sx}
�M���E0�iL��L^z9�d=��X��6F?+�-t�qD��o���1��qst�C���4>�j��<�����p��'B�H1'�����"�,�rȲ[��9g$4 ngV��ț��PCZ��s��z�:"{��r�YУN���K�j�Mݾ 6�1"�W*|A�ܝ�������3��T�N����Z%@o����������j�K`��{b�w?cqpk���ğˣ�\�5h�Go���lr`
�`xi����~�<��ʝ�q�H��S�m�%x�`#���Ĝ�Y�wV�z���&l���0�6�5�
�GR�eJ�ޏ(�L�jt�`�'�OQn�/�L<���Rʉ�_jҥdopnxc� �P���5�Pd�ㆇB�?u��������q��=��qH�����z�AdVp��T�����R�0�?aI�S�Ń��S,iϞn�����[3g�I��d#�����H��F1	������Ez�m��Q=��2�5���4}7ů�u��~�Ħٔ�qĦ��}'�݌w��
�q�S�'�U�P�����Vg'��p.��<4ׄ !���y��� ��
œ_A6E�>�P#~��iO'���Ay��n�)�	EE�t�:�����bȈ��R�Xh���Y�ǚ��i���TT�"�3.,M�DI� ����f?nƥ��R���I�O�&�t6����h�\,����*��?��4�BARA�1&�B��ӯ^YH��^���V{Q(� ?ٞ�h21vXԤ�gGy��v�w��t�c�'MxW	#���Fe��,���L����+.����qҧQ�A&]izN�!�M�R���ܜ���_��>�|;+j���&����>�D�΋��`C�$�՗�z�
��jf���l@�e��f��^�47֨eq���h$����o��X6�Or�	�S$϶���f���ӧ�i�e��ļ;��Ɇכ�~{�3�j�_��qNw~����0���/�r�X8C�X&n�A����Y���|����H��ajp�4��#�:���:]W�L�����})�JuV��w���JJ���z�NY/�#�N�ǐ�����IF���b���t����5��wMڭG���f#�6bf1[�\����s��CA6J�܃����S�J�v�ȳ��e�|'��b ���j�D����ks݉�X���%��b�[i�!.C	��A�����߷�Q����B�| �s������=���\zS����� ����2��d�H��FQL����û��Dȉ��l����^�Ǭv��XL��U�1@�+�:��+d�*n�,_��5�J��[s�!�O:�7҅T�
��R�eO$�\���+�x}鮉[D	`z�0� �Kd��c: +��W����봌���mѲ���B>�UP�n+�}ժ*-r'��"�i��:6;�b�����`���ۑ�+_��O+����e?��Q=��q�6]��m/�=�>Z�o^����p�e�ҞMӃ9�N�״�b�jL/���������
��v tn �]��X�.[��s�m����8��J|�E&��׼O/��{�Q1p3JڌP~Z	���5P�v]��V=�����������f�Km"��@)��CrN9�wQ�U���P4Q���N{I��Kɥ�`�D9B�,���;�ҝD �ײ�:)�,�(��{@�UY����[_��I� ���-�K�m� Px�67����9$>��8">P&~	J��u�E\�)m�!�(�@��Q2Z!��3NT~��cOIDl���z�vx����7����gd6�8���AF�����V
TBy((�qn��j����(!�p^`�(rA�1Ԡ6��������9���HM��[4M�v0_�Ae�5�<ks�_��x�N�qy<���`���l���_k�V�z��&(A�oY�Tf�%r*Y����}�[��l���Z�� �;��P\=Aj��=vd�
�c��wYz%Zj|==e@�k䤸��8�Y�Q,i�R)��z:�\$����@�m
��R��R�7������*A���JfWufE	4�K�ؒ<���ʎ��-.�p{zd]�]GgtUW0�"7�Jm�'�������0��T�f=Gte��!2�tOUP���g��_��E�#��q�D�r��ϣ�����y^z/�sq�OJ�F�l+�^*�P��������/��D���������vXۍz����|\�F��p�S �2��(�K�(d��ܟO�����b�HL��&8'�#	m��.r@��a��&E�^9�fa��`O�/������Q��P�M�X@���v�X0_U�\�<��E �Ҧ4v�C���dӨ1rʣ���ل�p���n����.�^xRB��T<o��ͤ�J�/��y�c?����$H��+����PY�:xJ�p:,2��S���T�_)���H�c�؛R{^�6�� �FbU�����Z�W�&f��$Z?ԫ? ����<I��_ɞV�/�z�``����b�0����Z�Hƽ��:��IOh�B:YLҭ��3����l�!�Ϯ>�?�ӊGbI��)#��$ł���牦s�7�܍d��*��{Y����!c=�e;�F���<�<��y,��������*ĕ�f(��f��c�qN�������(�U�j�K Waڑ��ɖ8x��5�[ܒш��$Q&p�
}ҌD�����R�\��)��?�3@�A�����?�S���}-0Ǘ$-�3Xɪ���ay��"�L�z�~�{���8Ӛ��P '�-�q�W`1������JR�kE<U2�� �G<�+I\D�����w3��-�U���'%J���'�K�R���z-��7�@U�p�`��,w"'����<����c�Z'����LWB�O<HO���������پ����Z��C\�a�ٵ_)MS� �	�.����$�٥u �L��`��F+m
�6{}��w�4�Y���!�����^m,j%�bC�v�E�ǘi0���A��4]�K�:�-g%�����(|��b�;7�ʁ�
��,l��z%a����{1�-axg��P�Ug��#�;���HK��JZ0T7E_���yh>��.���~��@�x?�U�i�����Ч�%)j"�3	i3Չ�T�it\��e rEZ�Pi�%��*���b`��ҴH_3���7k3����.H�<��%=��)���Wz��q�NJ&"�-�Q�!��JA	��U(�q��|YpI�]�
��i!}�>�M뭗��M���Ԣ.sT#�v%�/���Eq��2��!6h��6oà�����e�i'��a�p9t�.�1�p����VqMp<k�k������WX�g�"ޓ�w 2�ĭv�^B#W�\u��D��.2������U<��^�x!=j�*2���J�K��G�YΤ�V�/,�D��EjJ.o����_��*U_���������O��;3z|�@������;�5�������Kb�x���;HT���f��T�*��˪��ZGբѣ�FZ��#/:�޾|J�1)n��9���sg����xk�7���	(w�M�Je��#5�7��;I��v7z�/�F�ǧ?.�>��/9S�=�n^��P���5挽-���W9��r���㴖\��-���w<�6F�Gm°�ѻ�Emi��&�'34!q���@L�I�ڇ'�w�!62����u���/����y0�`�hI��u{�T�lV��7`4�L]k^R�Y������h���8�Q�+)��S�G�t�����E>T�a�'����W[��L �����<���f8�-O�Q���5�P�&��Jf���p�f�\���^G�y��7�|��Lk�=&��+��b��A|��dr}BVTV�:h��o�@=L�Z�%����9vZ�0��fN0����A��tfs�)+����@ځ��@����.\0C�*���.O�(Ĝ��� �������[�-��L7տ���A���8����Q<�R�����Y���n�_�,>��=��r?a�C�ߨ*[n8PI3~K� 3�b��淇���~A�o���o.H��R���>Ǖ�/�8�+����d���D]6�N%�������)��լ\��M<�hN����=4u�m�`����;;��i��e*v�	�e������4؀Ϝ�_�ȿ����Ԓ�@ ��MA��Q�V�e7���t+\z�V|�a"=ͯF?�5��ݠ6}Z��;/��6�x�V���.�\���g���t��hΛ���x����Y6]���$6pho�`��P�NC3��":��$/�}$ n�ϛR`x��`�t��z�(�035OE�CBo߾����2�&D��h���N;gې��������v[�&�A���N�� �׻N�'�����};ܳ6��Z"���}y�����q���1jlv7���K����#�9�.���O��u��P>V�]���s"��߸�å�M�N�����w?U�E!ɯ��,nG{�r�#_�M���C��k�`.�W�'ņ�i%v�{4�{g�Lz��m�oJ�#������0���B��Xy����ě��rϺ�ȭv����=h��C��U�j�)��g�zޭG�Ӄ�P�(�֏˱���Y����rG�_#,�,�Dv+��C()�[�S�7�G����c������h��\� c,�Ro�цF4��q>{�F�]�)�By� n�r��[��Ļ/T)�5�ԗ�zԒ�p����j\��j��'�ʻ�[}��c.�>֘�����w7}�\sk"�۷����!L��\bsj�U�+}{��:pρ��u�Vkpn%��X����-���mI�Ǧ2F w�"����&���Y���$3�xZC�{$�F*D@���NrmJ�3M�;{+�R株�����k�P�++��be�I�~u�OX�ʭH���RX�eq=����yH�8�F��*^\��T`�p�"�B3�}���b�W&�n��0,���<2�-\l����@ç|Ib��˝�	��/%�h��yǻì����
�>(\!$�zv��R�N|ktp���_��P�qFS?�rm�����ݯ�A��aF %��F=� �cú����7��R���1D=C�Tr|M�"��b�[HtV7���,~�O��*�S�cXuhe�]�h+���}w��΋Ј�gt^UI&`ӛ�	J&omdkb�~B��W�gЪ-��u�t9�~�7�sfJ2�0<t���U�hTd,���{`u�d�J��R�U��Ȱ<�Wɴ\r7����N�K��6T���C����W�����&g�:஫��`U�䪷j*��@�N��^Օ>!��.^X
��U��A+r��,&9!=�h`�)�o�g^�{m]��DUX����F�ګF�Z�xXg�pykl�O9���)��q6���r��,Π�B���ߢ��\>����	r�ƺϊ����3Xwd��j(��AY�h�}�e�j�RTXԼ����_5�3E�Z��;�k��rg�U!ц�Ɛ�2ψ�NA���2�cS{�����c, x�᙭�~�	s1�oɆS���vIu�L"�<+���`be:���M�����C�wS���PE����#�-6c_��:��U�+���h�nk[E�����x5�e�i����"]C��ߔu��^q?��֔S&Pqi}ֱ3�M1��r��ޱؾ��[�l5�b60@�y5ROTޥ%,�4�a'�����p"ox���yb6@�.���?�g#���ۿ��]�@�C��'_�̚�������L�ǁ�9��Ɯ��������"���&��	�Y�l/��B]����
l!k��p m���z�j��>ɸ�����-��ؤ"����<P����6�CbHø���m��-��e�]~W�� ��dA��� 0���9ŗݓ��K")N)�u?`���X�sW�#�U���ӺG)�ek#o�]1�(Or��r2:�	�],�n�a�Kڏ%I��L�Sa,J3��C6RY��[eU����ʩpĵ�z�@���Q�#����͈|dt%)�p/���_-�<�A� B[����e��-��W���!��t��B�1����˄��j4�;�,li�/�l#1%Ĵ������T���^m���y��)��^߇!�.\r��\u͎��iP�����'����)�����j���/^T��p=���/��[k����Z���ƕ�<<oTo�6��1��Ro/IlLa�x6|�j�<S2i���OtPΙ�*}����G""����f�"��xR=@���_�Mk��p1�Ń3�[� �M¹Q/������������/yd�����:X��o�R&n��Ff<GK�a�UY�Wϊ��2V	gr>��Ґ�Zr�����rH�+�=��(�h�|��繏�ʸ�o�E��5M��N\^:���3���*o/��Mw!$r>��E��ٔ��597�$��Vk�ǌP�at�`�v�y'x�P+bwQ�d>eaG�2b�� ��K��#{�R��J�j,��]F�;��Ös�	��l���s����-�[ï�շ�`[`O�^=��G%�?R,�ﱛ�wg�O�A��L3h�b��L"+����9�k�'h��P���ƙ	��V�+��Z�㛖{���%7��*�6�ᜩ�Q쵻�:�g�B�Qמ�K��~Iߔ��L_
���Q����&`ؗ�P�zC�nk�H��^�~έ�}$}r�1�;�֜�F����ֱ��r��׵�s>��:��w��q�oz?��rV�q�Ě������ D�0��8�u�:��g��H��>�Vs��t�6�,����k^�;(�>�'�=�Tiep��o�QFj�;�q�%I+<5�x���0�R�ؾ��}��S:2������ޣ��n�3Q^Mv��^�#
f��i&�KCGK�X�y���<�b��%i�������.��=��Q�����#�U`��5'����cϟ!�k��C�c\��?�&���l�]L��� �_�q��nU�o!k���Oݞ8��<_��4�}%���q��9>R����А��DJ�Gt[������U���)L�sY$
J��E�_��:n%�5�6v��`���"�|%���=���svtc��a��s{��#�ˤ�v��g8���{����lE_V�T�9�dLV���0��7���2ð�Y�.4)O.��1��{��@�HÌ�М�b�J׉6
���7�0�H��
�$����<ˇ!^wφ@�N���k��iu���|s�D�~Yt�>�^��\����,=8R�%oo�1��>�:q�뻣9vI,��)����N�<p���>�~�_��Ym˜�p�:�jX�Ws2�8B(��=�raE@�w�E��T�+!] �+j��_ʫ��{&��p,�Eb�m��$ǿ����i��:Ƥ\��c�sD;�S 85Q���rB�z."hP���]r��>Un@���>�DR� ���b��)���M�-�G$	7����bs�Źս�۶���//[YH��Vd�b���Κ`�Div7������UӠCc`�.�E*�?J�.[��@�N`2G`�D�/W� Wd�e�|ɷ��9�R�U���yfy��㉹��⒲<$nf��(Pul�oH��<�+�fP���yN��3����cTꅂ����l����[�m�L�l�w͸�O{�،p~>�� d�����Mـ@�%���b��vq����O.��C���@A�H��f�ľ]DK��#�O�Ձ<Q��.���tՈ���w��b��|�}��	�
\�jVG�,&-3WS�B�:%%�M$��� ھ0|PoY�L�+- �k�f��f��:]��I�]����[0�,D	8�8��sU&I��P��s����69��F�,p�`|��pP�:DѦ����4���u��j��+�|Y�&�
��MՒe"�Q�v�Bx�̟j�a�c�]�e�w�����5��qy���+EXv��=�,J������������b�"�#�S_�f��0�IE���T�'����Mk"���t��^����5*���'yF�.�Q ~)�H��,ӆ5Xé95�&w��@�6Ǫ�'�77g�d���'�!��\O��k�')6���J���>
��>ic*_��Ѽ/�r�?E)�t��B�-��-	-i1s��>�K�2p�M1�b�>)(����ƨ6���1:<C��^��d���b	�[��X��=��0K>CVC�����< 4�=�a��w�pR�v+k�T���ؼ�
�\FrRiJ�����]����N}����
�b����J�)�!�������7�۽�UP^8�h�ϼ6�P͊mO�{��Q��U���1p�lX�h<�Ue���!T���a��7���:״z�#(̯�MW��׭�ِ�6%����	l+8Ɏ�&����Yiv��� �9,�o�/��s2v��\I�K��w�]
�L��|g� ���v ��ۙ�a�KT��!��~Z�m8����_����o�]GS�۾&����'���V�,hp��N�z�o2��������E�\�C��h�*�?����zI��ܓY�BZ�,�j�WO\�?���Wz�5+p�_+�*c
��9��ք܂H��є�T���$���y�����?���=�lH�"ʫ���H#�p���9f����'^/��7� ����[���+S�������u��A��9c�w������l�Ȉ�x��	����GMyj�f݀8�ڞn��ߜE��+�V�y[S��rgj��3i��/F.�pb@�3�,6׶�Q�d���]��k��(\�#�5��h��Bb��o��5-i+ͩ��:���aG� ��b|�xƁ-���ݡR@��Q�X[d����W;
�2U�Q�x��o��7%!V���<�)xZ�z]@�tF����\l&,��&�4�������~�h������ݤx��s�����?�&9Q0wx�t�8/uTT0�p.R�AS��A ��ȓ���i'�-�`������t|(��]N�#!ؓ+4���*�E��Q:�-k�X��1�+ڃ���S��p�B x�&د���>�O4�$ꡃ��&<�Qu�/dul}Tb8�塭'�Π�~���?�%� �5S�3��jv��I�Wn�5B���������y������R���˗�܍s�UKf	�v<R
����Ԋ?��O�Kh 5̿s#i]/�q��*�@�3�|��Kc/M=����~ȌQB�T"����N���7�r[�ü�O��o�}>��-K<�Kk�&@Օ��8s+q�*�oZ��C�����m2Sx({��]�e�#�gH����>��uU��3w�1NGP0�)L�e�k�g�F�S��(����t6t���ˏ�J'K��M[���1Ǹ�TA^}��yJ<�`�G��_}���L���Աo�,�ۍ�@�K�-�{���f��7�/�h�Go
?=�����L���C�Ҟǁ�'y4y�{��}���"Z�wTF��Dq��$@5��]�2�F�Y�O�UM.i��wG�!4'��!H�����׉��!ol��}G�ߔ{֨@	�P�hR������y��h����w��9:��b��f��|O�b_�W�HG�а��jcr�צ�N"�����D8��[���H~3��f���;�,b��΍F3�#u^�#�K��E�L�Ѧ+���f�@pm�-�j�˔����3.cU:$�{��C��ni����Ǭ�@���I�yJl�`9��q��3&j�#�����;�yY��+.�?��5�بݒ���xd+���G�3,�a�,W�	�Q���֕�V�Y�2:J��1)x�^�Z���9R�$������qH��=�D�8�;ј5�\���T�҈�����'���J��t6�Y�����8�3�����z���1���"�[/k�$YKv�s��>�[b�WÐJx2������p�nβ��<q�����T�	�/G�ٍ��TXăyE$h���'
m�dJ�f$��M�H<sx]�c	��m�D��(��H��� H�����=E灡{�N��`Փ(]D���������/fzA���h<����v��M�@G'յ��hV4�S׸�TI$�O�(^�o��2����Oz�p>(��Y��Nl)/�����&�[O��Rd����ģm�H�D2G��s��1isf�P����6���2�B�W���0�I��{����C��ܷ�U�����L�*�g�A�/0�1e�F�,�onG�IG[7+�ך�(z1��%�����b���^XQɿ`��h�88E�dt��Q�eA<��r]��0��p�H8Z/h�4��$!�6j�y-��&,O��釡A 6RYmd���OGO�̶�`��!$�o��IAn#y^�kn�Mʚ@�B��.Ty�PlɆj��r����݀~I�8�Լ�\lGP�%�ʉ2q�1��3�7"�E���'����:ȳ1��^�	zwo��?T����f�٧�5�g������ԣ�����+�P���M�[J��rk+਄��d8��)�"���x��.��阕Dv��6�J+��ʄ�^P�"��ʢ7��w������
����-��ۦ�uN���C��B���AY��bq"C}|�qO��%��ɓ[�oھŮE��E5X���`�{�VGu��SQ ��������*�x���YP����U,���Z�	#�&��;>�ꪧ,�'O����c�^�"���"�y��u���oe�M_@�b��tOR�,I��&��K�g_��|C� ��A�����	���r��P��ć�k��W�#KF�F�W���UYp��n�aDBo���a�
�y�h���3�D�!�o}d�Ʃ�����*vѿ�ψ��'���P�khi晞M;F`s;���)A
R-B�O}l�k�-a��X)H�¥>�W3�J.k������)ւ�5��Z9p��~A��K�
9�R:�JF]�dV o�I_(��6H�ƫ�<0Ez��cٮ��Ԉ��W	*�dt(�fP��,���ȕ������E�������n��(J}�q�Q:���7�'�v,|�N�1�J��TgA���Xpm�Jl�!;N�������c2���(�a�5@��" �o���Jث�YEȦo�c�^1�t����5�G�|}�$�A��O�Ҝ��������tg�]���r���7�{��o	_�n8�Lm�Bb]�q�����7���@�P�ޢn�g0�"���S��]٭Z��y�[2Z�sr�˛�J����,ĆIw�5��gɟ.̝o+)��F����F��c���e�NB��S��C��8��9IB[��9�#�`I'�K�N�p��t�q|�4�� 7��0C��`Ԭ�~5��g������/?� O�Ǝ=i�	�s��lY��s�0�E�h_)�
�-4�M��,����T��3tA��1v}����*�g�t����c���"��_p�7h�Q{������;(��Ɗ�!���:����t�ĩ��;��)�P�4h7g��tV�H��4څ��ø^�lRaMO�ـ�R�z}�\�n)�����2�z�˕%5຾�]j:�"�M��d��we���ۍ�/���M���q�yz,�9��ݍrm��r�O�(��[����UrY�\�T[oޖ�q/y��W	M�>�0�r����8�K"ꂲ#��ʶ�����T��ni�����h~��蒛�w&��ŕhC t4�y�ޑ�D�_,a�[��6�loD`g=P:�WK�wTr't(]x'����֯�h�
�5�aT����Q$Ȯ9��w9�X�ќ���
�F�T� ��}BI���-�o;��eYZ2�n�̺Y���3�dC�����_R�x�3H���&��d~�T[Эa�΄�m�����*��%,yl2�:��	��G�t�p��!��a:��T��@��0!<p�"s����@�Fe����4����Jg<(��Hm��Vn׉
�}�8�Ǡ�� cH�>?��\)KS|{�.6�C�I�P�ݳa��i~���n8b�n����H'�ё�+-	�H�<f�&��m�o5HB:����{`ބΓ+o�q�s[���Ev1C���)�/�u�Œ��k���w?���)7�ԯ�n� #l�?�1`þB�,B���{Q�G�Kf."�]���V�A{��.ӆ���e��DT��Џ K>�G�z����|����h<��(���L�2�H��������� +HJ��Ԟ�U�� 픠�,�H�m�8v���Pe��C�v�3������� �jȗN/v����A�`d z���z����Es�-����Nv
��7���|�y�:c~�΅�
��_������	frP��i�<����SKi9Ԯ	��֚�3[1���}`����cd�!2sj l���W{�u4����_�L��؇.���"Dh�"r���O�qޙT�b�D��D��$��6h�:h� �Z�e1BC�2+��oF��+�@|�U��/���I��)���zS�v	�g�LA�H�~i-AXs��䴥���cbH���h���<�z�&ޕ?���qL�P��z9�9�k��ƹ��4'��Y:��ӡrQÿdX]�nj#<��d�~ou��p��ĪM�?ڒ~��خ. b��O-�>D1ʗ��Hb�k�Bu{ HɗH�u����(b�N�N0@����ST��ƭ�a��q��`)��7��`�/�� �S�Nm��2�/��!�,+U��A�}�E��}�(� �N� �#��^]q$��|<-�,�G#*�xD`�8r��@.�]I���LK���mh
�"�u4�YQ��Zӑ�@��,�⪾��a�߃�~W��vj����J,+a�9� ����|G!˳0����X:J8�č����@t[�g9��7G�FM��//�
I]����vR�2*Ε/���d�������� [��]l�n�H3��R1x�C`��Z��X������Pk˞"�)rk0!�N�;���s�J�+0�Lx z��E��U��<R���̀ͮ��mO�k6��ū��[ē}���ֹ;D��d P/I�Au�Vj��)��6�������������@}VZ��p�O��NCB�:��V���$�J��w��"�n`������i[Z�G\����'��{���Z��"�J/�4��G$Ť���$�����}��D�G@Ź��z��±��0�|@��vp>�jk�/�j��x���R�o��&Z� b~�x���4W�l�Ų��^|_�5�n�B�*�}ā��G�N��;�������ӑ�c�-+#VX�`$�O	���y�J�7����I"��Ѽ�:��y�%���%L��A�"�m �/�*��M:��]����Eau��]��0Wy�{m��)!���$���H��L�
�7jIyx(\fzx{���6д��Ye=_�Z#��;A�\�1��\=G=\��_*)Q�?+I�)t/NxX��{�� �\���� /�!��U�c�/#s��=����9���gл�2��r%
 �g�]ux(P�����GU�j˃3w���T�nj�K�MA����У\���CR��I�8��yt�H�$J�NmfjX�P�/�{�b�X��Hl���������׶%��4�`D�b�8�M5Aڪ5׿a�Jf�o+w֟��"��s I��A���J����*�swX�hD���4x�Z�R1���0���y[�}�Q�dg8�hf�E����͜<�s����>(Ӕ�#�r�=�'��ᡋ��T��I�đF��*_X�<I�R�R�7�D:e��]bK�4:(��u�Ҹ�G�OdY-�7��dC=:N'siz�+�9�g�Ϩ�3�舖J98�}�]��Lgm�Ѝ�?>c�_����'�Ҧ���?�B'�UD�jvy��.o���I�?��VD!i�GJ���1L{$	�.�[�\��C�Z��bJ��D,��W� ]�2��|�Vn��`X�D�8�q��|�^�^؇�fT���5�SK�$�tq���A����V����}�J�����Hǀ?_��̧Q�#y�t��Q-�b�l�e���fP��orv?�f"Ό��yE��_��F��Mq� ��ɼL�W�.i���C=�`�fT�m�"w�6���^�����F.Oӥ�|q$T��}�p1�4xZ?.�I( �3N�K��������_�,����"F�,���H�@���̜hFW������Ř�V��&S�")z�3v��rq?��
4мo�'d$�Y6Y�9)�q����(;7�����bX��w�NBd�g�m�bGCr'
9�2�;�AP��kq��#�􄖹��C�Ew5�F`�Jז��1�P.�,���%�������&��Je��j���ULwד{�ua�.
?����������6��)�;:��}tSBf�~��L�d�.���������NY����V`jRC6�ɣa���(�q����)C��7ᐈL}uo�V��;����D�߻f�X�}R�&�j�1E4"�3bm�R��E�W?\��i�u>�[������Aaihw7�T���,�v�A J�*��	���xQ���F��%�Õ5N���g��.���	�,<]&�4
F�9�o�#dT�EZ�(�0���,<g�O�d,�U#�xU��rOk�������I{��VG���J��O��f���Z��X�n2 Z��K�$ �*��fl��lx��l���I�~��EػRѭ	S��7u�L�Xz�8�����3_p��y�jJ�սk]FnٍmW�d��o�����Ӎ���tJ�m�>���x�M�8�L'.�������$���'�eA��]�[7 -b��$N���@e�J�v@U�P����hO��
 FN��Iv��A�
�2��`Y�bƔv^���kRP��x�c��bj♋Q�n[������e��z`�ˢ������Q7��� �o�Pƿ��@O�y`O!�#meA��/��T\%�KE�J#@`o
0m��U��"�Z�nHO֢f��fU��J(Wa�rq�5y�f��|w])QdD�#�$p	��2s/�pŰ����#Ƹ?NK�p� ����'q��Jf}
���`0r��[�H~%�W�lbԲ������9t_P@��K~x��=�,��j��z�Ogw�[�q)r�ٿH/Er$�5ݤ]�zm�Z��-]l��9���mW���=�z�l�#q�� ��8��"q������0�rӬ�T+�x�X�觱�����'�4�a�bҬ������."c�~�P�r��#�R������+�/����_�r���밎��ɓ�4 ���:$�&])��{�:YՑO����6�*�tX]�r��P�aQX�R�3t�ۉ�����{��a�|DV���n_�mx<6�cPז��;�#h�GŒ��е����+X
˖����E�m�RpO����o�E^������?#��A�~����n=�i��[�4gTB�;�V0�?7��4��C#��d���Ka�n����y�&T�U��}�|��Z�'�)H��1 ��3���CyǤkOU��r�������lsD-=q�O��W}��Y돔�ZV�IG�B��1]�~�j��:yWo�� �r^��|��)����f��|d�����X�뀹��U֒1b�s�k�GB�!�C�0�v�Z���}D���^��~���9���{�ʍ:��ٰ7*���`=TZy���x�I"e�.�X	��[�`v��-��L�o�E��s�.q�`���A)��g�!�o�����A�eCT�y��?�k�r�|hT^�C�1�O���H+(���*0�u��%y�P�.^4+�К��&2࣌�;mh�_To��9θo��EӇ�P���z�#�����CM�*�x��2s[?�Z���M�3���Ԍ���s�f,�\h�����QG�J%�
�� ��wk1@i1�Ll���k�3`"�� ��]3l����Bv�C�"��_�)}u^3Ѣ��'F�,�����:ж�0�)h�{bٯ��K�0��)�X���1�&�7X~�i ﯹ�����ʸ0���Ij���d���MCf^@�k���� ]�`���O o�o�?@���$LQ����yS]]@  	as�h����</h��DV!�G{d� >�#�/V^e�+��x���`4"5=�^q4L��j��#a[B�SCP�#vB0_	�1ej5%��ɸ��2�1fIS�w)5Bj��f*����\Z**�G�C<��>�4�ὲ����?>���D����Di/�-E�B4�i���[���a��K��_�Ȧ��?���x崼v�6~�H��ˢw|� F���ɠ�IN`6EW�k:��3�	b�-��Рtû$�W�ě�D�S������d4����_]�P���q�s��F$\��F��N|5V��\Ve����p�>
�ӞBy��d; ����2cr\��N
z��V�	���.����~u���(5�YK��c��ġ�q��'� �<���i���cw��m�?�H@��|��-�k��5��+���A��_Q�U�Y��w��Yl� �wQ��V����5� =���"T�I���+����LQ̧kAsb�P���Z��;>�5;���5�ɗ�'�Д��(�� E�&�@[�@��
,�(@/�#� �ӹ��I���?	۩ϣ��)����K�	h���o�#���/�iP� 4ؠ�v���AМk�zM�ÊD���梐�Dn&I�ދ��$P��L'�zaQ���$7�&�!����l�*�!3`��R+�:���W����1��Cf�{�Hܑ���7M~�y�7�h�Q��͟��7���B	k����8O@s�)�o�YF�{ģX 7�^?Ҳ��!�~��CuE�b�F_�V���w�p�a|V����q-����#��+�TE�7���D_�?���ױ��w��{+�[��ay�VZl��(k� ]W�ݔs��W����};g8���_v����g��^��Mی{Ā{mՖ�sE�2���M�[8_��;�]����O������\�&44�ZH��{����Jl�s�b&�u�K?�%��b� Fi�;=��I%GbO�܌G튵M���G�L�3@�)�'�?8�������'M��U�a�������G��!'Y�t��mڎ%_/�(�f�iC=Ü>�U�ml�6�,t! t�M;�V秣��b���9 �9���l
ިK��p�P�X���&�F?����	u���m�i������6�}25im_|�?���n�P!���%W.cUD���G&���A\LNݳ�$=X���1�J��'M-}�kC^�d<�#$\M6�ƫ]���Z��.�X�{<>�e�������(''�Z�T;"�e���tpBdaF|˽���ׂW���㗸[�ت�+7�ؾ}�����E�������/
�.��/��]Z oF�ɏ�FS��D35ߩ��a�"�����R�����.���(y�ok�<2�LW�t�0+A>U��*���L�p��Y��^�<2?᫟�q�OG_� ��7-ZR�z�z�����WڽEV���/�C��0ߗ���@K�O+i��W`�at��@���YD�䎀_�q۽5o�K8Ξ��\�63l�t���z&�47΁���<b�ߢ���hOf�7ޟ7��F۽[?tl�o;J�O��8v �������<�[�M�ld�V�;�c���$�2w�zߠ��F�ëy�d_Y9�^9�<�:N�.�QC�V|	�"�Uvה'�z���T����1jV^���h�������lb:g���P�d����IO?:"�2����(K< 46I@�]�8*�h����\�s�h�3�M���d#�x�֣��l 	��8�Z~��,���`��zU�w���x�ج7>��x��ʭf���|��tP0������|
30oʣԠ���S'u�Vda�&U�������
�, 1(�Lv�6MK C,-Wf*�@�B�_�����R�ǃC�������A��*�F �XD}b�A� z�;�}��E@�uk���*�V��~��	,wVB�z%�&v��Hv�z�0U�d_')n�d<VT��#���E�V���g�^�)�Btʟ؂Um���L�Y8�����-<;̪Y��\V�9K-���K�m����A3xa3r�&���u?�5n��U�ɘ��)��$J)_׋.���x�T�[ؘӈ��$	����SQ(�
 N��߭�:M��膕W)o(~���n�_Y3gw7k�{�����Z2Vk��
 �VԵC�i^��r9h�LǢ�tQ�WX�-�P�~�/�A�;��IQ�)���u�V;�>�9 6�q������ȡm��6≛�D9�a1a����{It��+���`h���F���w���F�#�a�4hf�$2����eT�Z'�wY#x��)<!�~�&(�i�J��=�kUI�F��ڇd�L޼b`�����ԢTG���4����W��T�Gݠ��25����;H�va�&Jq���h��9��;�i#8nJ3Li�_�t�+D���X
H [��n�����������
hh�>�L+���,6O�f�t�'���*3*rn�M�����½�<���QH���Qr!�g�F���*��޴dV�E�i,��>e12o��xMb8��	�#�&����������Sy������	M���4X����
"&��m��&@���o�`ꭎa�.����
��B˧���h���eL� �e-v"�:��n�x3@��=g}���H�V��d�b��m9��)&c#�|].��/m@1X��OraiGO r��~��"{�0�_����~!m��5���a�s�j��V(�A�Bn��t�����.	��ѐ�{xR�-K$��NON���bx/&եĀ~�l?��V�	 ����{ "�{Cf�k2�L��+}����Ů���R��QV��44K3��p�%CmD��f8D�Ha�?�D��s��O�	�'S�*�@��㒛�Lt&g���&��#�W�����;^9ek�������X��.��q�����CH�,؞a�>��aC5�"=��Zĺ����F�Ǹu`	��+��jD�:1�9UHbn��D����.��HD��4��cZ>lB��/���ٛ��	���g��'!/��<\	�����¬�?\��тQ�Z`J�;t���^��|�4� ���k@��	U��̫�@FG�K�y�B�
��[�L�) �L�7yy�@Ўx�?�:�SW˻8���<�ɯ�%��-�V��7�6�6U5��AaR�i�����i��-zr"���6A�?2��r�nى���V�mO��W"�v�5S(i���8	����c��q!����b��^C<)~Y��q��eb���P/���\J���\	Eޤ�70����-�B�0hL����2$1��ק;��H��x�[��c�Z��K�܅��[|�'Ɵ��oG��:������;�j�z�.kHN�ڠD
4�f�35�d�7��p�����M$�L|��N�f�>1���voW�&�B��n�{��;�k�Rh)�F4�%A�X9h)Ba���dw.�vA%C�W�X�)���֙W�%̬"�B�A���o�x���+��8J�ʼ�R���[*U<��V�D�/A������‍�iø]����W�BS��`Q[�@1��_Ϭ��k�;*�W����yK�V�}����]Zג�DK�\>ѣ�P��<iN�����Q�]1�b�c����i���R��].6|?��Ҷ8�r籹/�Qe�(��l��@m���6�(<�|��ی�O�bJ����Mf���1N��l^4M-�<�q舧h?J����10��p�@j%6[f�󥎁ľԡ=~2=�6[m#b3����!�����v��9��ȟގ�@?=/�s,^�rf���P��1���:	�V�sVϕ��{���������>�yN+����4�����*y%-��)d壟hb���L3�E��r|�*��
1<9��Ǵ2�b����볈EeE�gC2�(}:���F��爓����,zȅ^d�o���$�0�p��Â� re����������aU��t�(�$��h�>�� s��y!���������*�}�N����t[-8����ǽ�<2�3ӷ	0�X���l�y?�/w����������G;Y��#w:סd���¿dM�K�|9 ��+3
�H�O��:�>��]��g1�c5Bv~�%��}�GW>�ڸ��ty_ �[T�#��c:��JL��~\�ל�Y@K� ���T;зi�l��.|F#:�d�4|�Z�+\@`�z�Y�H��\��F��i�e!���n�>�g&�q ��?�i>�d����z��ɓ�w���5P_F��[1�SF���������1�-�&��K=���e�{�[����~(���	Mx|�eӬ��Ƞ�a��q�_>\���$l��z�~�}�
�����a %ۅA�;����1�`ػ�����BI�1\ŧ�0󁗦$njoT%B0&i���F�%X#�ʃf��%j��Iq�	q'i���$�'	p�������-�8�CO����lۣ�xp���?V��$��!��'1�_NzvI��6��JkӸ��դ�����4�$*�&��&���KՂ�2o���n����6v��'��/��g�*�V��%�xܢ��<��+sQ	��R�N���f`�u
�!��L!�Sn@p% ��W�"e|>Yx!�]�"H� ��m���[�6	�*�*ֹ��+ P$�)ٮ�����.v�~g�J��;�*�ĉv1`��p�iz��!m�V��VO�+QG�d��6���Yy�2���~ ��hdz�R}2.��?�uEt���A������s�.9J �S!����nd���?��bP�1�ڲC(^��ը}^�W��[f������So9�%��p5<V���#���X[@���/��Ax��GR7J��{%��i�n�ߏ�'��i;*S�z}t��h��-#$�pE�}N��}Me�)��� 0#*� 舁����W�\I��C��Vo�MŖER�oR���c��􌸎���!��s����u�����e��i{{�Z����m#
�*�I�F*�J�2��x�e�JY.^{S���U-�R�x<��ND��uE�+�����j�n4��Wv��/�k|~���\cS�G Q1QN�f�v��s{�f( �SM������66rxq!v�N����ʝE�:�z�Y���u|��d���2[��=iA�em%����!�<���.��!������v��"�]}���~ī��� D�Q_�+.f����|�s�u��Cjy�8�V�$�;�]�p�l�!#��a��T�V<_3;�������K%
2@�|�_�v�vϝ�.�&�(�zyqQ�W�j�{Bm�bz�J�ӯvH�r�K��4�|S4��S���lmt�r�Z���p �Vz,�s��8F@$Y�ן���aD�L�58��/&o��=Oօ�ڳ]� �;���u�*MD�pr���)QXE�pN5,_�{���l�+j���5���o��j���u�E�*=i,3�]�)�,�*,�Em|�)Ž< ��H�Ys8����oo��?`o����xC9��b;��0��=��'T��psc�y,����(��AK�g�Ǻ���E���?������"�ú�M|ː+�P`��7/BR�Voz���e��y�厩�j�W"�^�@ވ�÷K�=2Oe�Ob�%�<s:��\�>���d1�ڸ���+�D�t6���B��:E�H{���b���)/���DüIPϣ)3�.B�t�q�K�%ɡ�M۬S(�?��C)�%���~Ǹ�I���'�8���H�@M�Rs��~V�?2=����d���i�yJ} ��9RΡg�r7\�����j�Z��L�J��j�O��K���@ط=�W~c�u� \�����!�U1�ʶ1�Q �F����^���	�k��6�-�۔/�!�9e* ��q�����=��N�(�6��4�"8����;n�l��m�ճ��Ҝ��~,���[�K���ON��C/F�]�{c�F�Rbm ��v-Rn+�������{�⽷�b��?{������8	�{�GԬ���O��n�������K����f���d���\���`�7j��8d�P���`c���&�0�q��,�'	��� ��4���h	qG���~	+|tM�0l�ܰ,�����=/>��c�t(�oJ�{�ɭ���r#�5H\Ge���� ��f�h����^Hr��9�Fo��џ����f�d�KL�m��|\>�P��D ڴr?s��7�U�sGς ��������*���j1�%@���rF}�M�V��MT$x�xڵeX�5�3���8��B�2�ǷN5�`(��w�l@������ͬ�/q2��'2����廤��U~)	�Հ�,Rs��ZBH�::/�:�R͊�N �g��O���;�b�!4S�����F;*���R�G���F:��3��²}7!���ԡl[�poc�E���v��!=TP�����������mfmre�l�t>����@�FO�z`	�U&�|s�0��M����v� ����~Y�/B�qpM��vfJ S���L�)��u�.|Ls~:��dU�����ݜs�P/IH��Z�v]:�_���L_��d�B�) [�zcͫ7W�����u�Q'_��(m��\�.h[P�.f�p��O�'�x� �e5駏�gP0p@��I�V�t�ʝ�K&�b�mMƱ[S�ҽ�.j�������=c���u/��[�r�H�F݊8w�'��$.��J^��Γ�9��wn�8;8�`�s?��x����u�黳KE].x���aY�L�L���c@[8�)�y�g��!I|;5sܲJYM�P�9��bڋ� ��(2�������z��
���)~�����!����F{(:3�~�����ΪH�[N�X������bO��B�q~�荴�Q�T��\���U�#o���y�\���U����E�Eq��*�М�����Ⱬ�~���>�p�H���|�Kz��tTt<O����� ����AK�%�c�ZY@�[�'��;�Sa�(�$��>yGK��n�#��؀~���oc�]�y ��� /!D]�����[�x ]9����L����	m�3�A	�{���5"������ea~���FY�F��f�@�/��	s��ee?�+4˕\�B;��5�+#���ꪘ�֊����cvsG2����N�P{��2�����b@��r�W������Ahrgvqe'�:$�M�٫)q��͋���������w:�LC��F��� �!�B���A�H#�����K�������J��oq�8�>�B��@C'pK%u����t�y�e�ځT���.d���#e���ط%;=-�A�oN�o��Cr@���� ��2�	�/� ��	�-?Q�h��;F�X�b��$t@��W%	 �=�$y�����߈(#:��.%R��êu|���HA���Ѵ2S@���״��`��P�������&�T�b�|�Ӱ+��b$�[}
�S!D~%�,$�4x�SH ���_]�]Ք|l!g���Q�إ�tO�I�?�؛h��`����6f,�z�O�FLH�K���_;I�Z�7>��"h-�c�f�mY�I����e�!Io�7A���Djc���"�9�b}�9�}.�P����V�m'���$�v7Ȗ�ܫ,���o]l��ӀP����]b�����)�l�!��qCjʷ,���c:.6R�u�W�e6>xKɲ�J����^�JuBr�l�ՠ�_��p��`����!4�����t���N���"�Y����3mB�\���vI��Ǡ�z������l�S�\��Ja�ҽ_ogT�����i���5����ݫƤBqm�/�H�K��MXn%��B;�{���9<\�kc믮�Ͼz�3��,��=�m��w���8C�e)Yv������ԕ�ǵ+Do}�$��HC��ԑ����H��g&b�B���lW�2����7ŘN��.����ה Z�9h5�L���`HR� �g����5�ޫ���d��������^�����aِ�#OԎ��B(��c�� ��(��	_�
r���oo���DR�U�YHV�H:�w��f+��M�p�V�,yΓ��siϵ]�x���^�}Dj�R-�[����c���D�tn�&h'�~!o��TTr�� ӵx�?���[�|IBA�!���c�U��#�e;80�W�("M�t��� �-�У�-3k
٢�J/H��c�!O@Xy� ]ص@W_���/u�bO��G��=���Z�s�o�B��i[�d5�\�����=%��'�S!
�#WI��|i�*�ݦ.�� ضɼ��l��_��2?bpح����]�Ӛ<	�O�Bm[!,
�5��3Q�)�Ey�礧'��j�kCȟa��h ���)��ι��Oz?'��AUd�|��P+�S>�	�e�:w�Mwj͙�����r����!4
��҉3�+�~ώ�SF��)�$��g����2��Y�Yn��7�`�[����/y��9�����y�B����ד?Y��\U��[��r��>�b�p�'�Z
(�))ӄ$t�.ȡS�Fژ�׎0�P�a�bP�IV�_�b�l]����g:��0���?I\I��񦥛/,��1���Ϡ�p���kA4%�7�J\H�T-ҙ-�^k��^R_$m	'i<:����=��0��@4��v_0,�op��@pf�!���p���5��1!_��o>�f�&�Z[rM7L�&@�@	��u�{�֌~�*q 4�Oa9���S�J��w�42+ql˰`�ZT�?��;F`\���d�+�¹�*}G��Q<���P{�������3T���V~]�D
qw(�h�ْ�N|��#�����f_�<2hOs��O{�xI[�\O�9�̨ b��ض{4Ϙ��Fa���I�,D�N�
'r����	�_�9�gm;ǵ7I��=,�������VQ�{�/�ž�ײi6��/���3R��˶C��^��m�R��IW�8��oj_{P���j�n�][�	�N_�^�{�k�����\��xZ蹆�RV���g��>k���$�.Δ���2m���������Z)�E� ���loR��	m�6����v4��|;�����Sc�ٝ�2Ë����G�	�V�#�`?�qI<b���]��Y,4�Tl՝SY���������@VmJ�:���j��h��sBos⌍�4$2�ĈU��m�oH.�ϧ�Kd ��sB=�"�D��ٮ�y3cIܬ#lְ�~�8}�4*�i�*6j��hl�7Sʀ����)�A��!�(��L#��>\��m���6�iNS{,:�F�X|[U�	(�U���?�����J�{(,
?�vع��e�I%�e:�5�ָ�0a�K���k>e�e�ׂ8У�,<Ɣ�Y4&V���F�<r��z�#����A�Ye��L�R�'�9�vs�X�ɉ� D�A�����a�	���Ys�Tw�M"��7���D,t7eU��- f�_�@�,��5Ɉ_�w����x��Q1dɴ���U�v�_X�&�`��DȄ��e;���Х��r��:�Ł�B7��%W�Hf)�������=8ᄣ��b�Ħ�V\���G�1)�E�[]@��9m=?��:�,�������Cʟ��U�L�:.@���G��ݪc����d��v�qc1�E��&vó��H���E��<��G@������T	C�,���bZLj�%�	X�ޱ��쨇�L>�f��^˕�fjEΑ�1�r==(3AZȦ;��/��I���ԡ6P�٦�;�Z&p� r��eQ�wJ�ވ�8�*��֮���5&׋H���Jz���ߪ;='����*=v�ߐ�T�q-��@�hJb����� �xH���I��<i��h��@%� �f7���JS��vĄo�"=�%;��,ݔ��Lȟ)������
��Q3RW�H��'��P��˫gan�%La!h_daQۿE4�hz��6��Ck'�@� F�>U#>��EZF��,����.��o���G�]�lC��,�"�����S�/������f5V�;�d�,�8>��Ȟx�YE~fjE�a]f���j�a�t��|�\��P��ݨ��N*�KQV3��؄�����?����g�ñ.��L����#�-
��XeI��]a�X��r�E���S(�b9a=����U�q��������P�L�LN��{�N6_�gݠ2`E���_>V�,a�&�1׋m���5;z��.N�̟��x��)(��oN��2�}j~�[�ԋ�ƙyT�|
g%�2�I)�ͱ㫣=Mju^z�oYrO���$hѦ'O��S��>!���OUw��7��L����P]x"�!aVu%�-|7�) E���A�n|:�8U�|��xW�*è[4�cL�a!p�B;߇���y�DP��1���I�t���"���h�v(.p e���D���]��!�3,�X���-�O�`�`��N'%9}����!�^Hܠ��u�!;��ԷC��������q����T�l���򄺩����4U�f��-�C^��ե�W��C����h����)ϥ��k�4�	:n�$�쮕����sL��ie�+A[*J��l	딇 F�u���̣$-|t�~5��~�1�Ǳ����Fz���4��0��$ =�)�< 4�a~;�T��J�]�V�sj<�eõl5!!�1�~����B��y����&�;Ӈ�6��L�#���e�a�z��䖽�z9E	(�7c�� ���z�}��5���$k��+6�Ē�S�*���+�9�D'*_��d$/|X�ɔ��?|q �A2q�t���q�����!����%�t�q��VJx���x�tc�ckz�44��R;���+��Z��u��u��y����lI�4M��J���h�=O��[͐$iU����S�:D;3iHF�d�֙�Ua�`F19�4�
����e��U^�Nc1$Z|G5+A�;
�yVa�����ւ���~4@d��kB��-��baC����%V��x�I`nz�v�����Q��H�r1�K��&����D�t�6=ɢ3{�"8
7a�;�R��n��֡! G��E|Y��F�8'��s��H���f�{SYhɒ��(vu̯�����e�k��Nw9߄M��s}a�C��(t`��q�h�u�:�_< �����WV���e���ޘI6Voy���5��Y~7ԨG�D��;�~:0�by��4r�
��Ue8���������f��{�-c����xo�'�-�"�������j�_`��$w�@nA�PsX�|�����uz��S�������8S��};��~bl�|�PvF�٠	�v��j�G^i����{��܊�T@�Rb�5
��h�2x�:��ë!����F���02�hS�6�o�$��]�<@h瓬��|d�aia[���8�_�WV�r4��E����U{7��~W���,��