��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)��<�=�!ʞ�C�Z��yt�vF�;[Q����e��Y�7W�/��̆~\��"�N]�|-��z�f�}u�ٗ�+�+3���,�"Tv��6u�)��I~�<�'�Ӯb#+�{p��l����Q����%_ˑ	�Ͳ�t_,�o�Վ��sz��r3&F�i�[���۩jV>rCWTuג�U���� ӴFy��| ^�n��;��Z�|h�!���#����3�8ш(Yv��f g*�BO�e�����9����p�s�AtG��8���0�R�2�B��� �=Z��	V�~�W$�)� �VӃ�0z)/���O�7�5�&��F\9�������QB��֛��>~���~�ᨬ{֤8g�˫����He巁,(��c���R_o�7�����z���e�Y`g�����Q��k@ר����
�b�hw�![.�B �Vm���'�X��{D$=H�˷B�h�k�dr�_��|k�����|]��S_�@dO���X\/�����Y��¤��ȶ�����3��mb�/�*d/�S����[�oo9����{m@�٢>�E�I���]3�qě�u��@���	'��\9���>6��U+�շ>; |��3�Y`�q�$�ѻ�;�$�����_�T}�b�:X��җ$�k|��B�r!<{s��Y"Z��p��� �B�G(�2l�G���Yq��[?8s�!!��J�����٪E6�nM9�����3i�`��W��g�X�j��::��N�������\��G�l~�Kw�� �X*�ݸ !.�{�����i=y�����C����=���h��'ےkC�*ۺ���3'�������;ם�dCDM��'1�!�h�c+k)�פ��d�� (�l���ܒ m�-߮B=%������n�>�f%x ߼��	�A%Mf�=&*�7�
>WN�i�ͬ��՚Dkg�Z�죊 ���l���O~`(�vK��$��Qh���B����]�����Mj[Ѻ�,�*�����rRkt
�Xd��cI���kVeˀ�ί��n�d�E{���2iO��y��o���!��խ`ae�X�t��r���x_+z�r���s����n�zi7�T�0dW��)����ڧ���R�N	/�N�Eg����W��[�7�	�y�dW� 	<Ie[�km�'
_�r�m,Re�])nO\n���f,"����&�b��hO�sxp���S�'�A'N3\�c	F����4!�6��]�_I�rGy�{D�焲�А7�hi	�Ԡ�a6C4y�>6��@�}A�ĨQi?�*�r��� ��O��5Ϭ���x��=wI/&�Wx����fbi����qM�h�el3O���SD��i�[�h���j�5M4�PS��1�@q�pu�%%�����p8����W�E4�Z^��G�<M�{�q]���ݞ��O��.hڣ~J���\l?t�S�Z��drb`:�g�]!pf&4�B��Q�D1�ۍ�N��$ߏs��f��^�r�x�n�-��>Q����ULk�3��cfPG������ɢꂛ����~�(�Ej�M.$02M�ќ\Þ��t���IE��۩������a�܅�'���ѧʱ,�WivOO�[�%�PX��T�/?�T>��A�`�,2}M�x��U	���.yt鶥�#��G�k
v�mRQĤ�͠Hl�v���7�!o��
q���?���%rK��-d��&C�+f:�v(����"�Ok�|��3����q�l3M%X�s�5�Q��Q_m���������2a�XF��{��W�L�Jf9���jB��w��+�s���Z�]dq������Cԡ�dv՗S:�֤ad��C<���#��	 �>Fm>D��:����������!�F;pM%����P�sr�2���bf!����~c(�~L�/�&��_^��&	�^�H`F�(���oºk4_ ���\a|�5OT|��5�����@=���y�Ұq��)�g�vG�R�0�:+�{,Pch�7��з��ҺB�`ڧ���#�]�:�O)��:1T�,z���R�Jj2ͦ�G�	
>��hTђ�5mW��{����O�QOL�\QӹN��C|w�ø}�V�C�x|U��*y�r��]�X���^��Q���jg�^�KO�Rhw� ���Q�g��j��]��/:��1�ƞ��Wy����ea���/
���g����!:�f�G(�Ч�2��S7`�U������8xQK��U�C�qr��0��Q�m�!sT	�t9WCc���?<������B><x#���L� ��i�~,�.�#h9p��ʝ�M��5:U�)o�e��R���C����>/�����c��j	���.��7Z%��y'�|���(Y_��Nqi|�s��L����ɻ��z\��[��m���2�K�e
26%��j��Q���*��7A:�,�a%���.�=�Q� c~�3[� ���~��{�-�pܹ̲��4�/{��56>��/�G.��Ĥڻ<��쐻�Jg�2H��+�H�Lkֺ3}�����F;;�Z�b��;�3[T�_D1�B��Yj[�;2};��i�����SJR�{ɕ������d�8�kw*���LX�����^T���S�T����A%|+���QY���#���}��3��:x^`����L����Zs�T���5�:�����Vp)9P!�A<ܨƖR�rIp8��U�|���Ϥw�����z�Q�����r�ˬ��:�b�,�m��ü�=�����E%k����ѵj��d�M�km$���d��Zu`!yP���
�$c��u2\2�����H!��n�������W��[r����\xg6�*�ͷ��yVB�E���(���|񢄜����>C�_먕*��H7u�}��B�%�(�1��D��,�3d������w�P�suWz0E�G��R�h:��'�uG���R�6�hդ	��ݣ��\��D�_X� u+����2Q~����8%KZf�$U���a�gr�$�4 �!��2��� ��8�Rk�.�w�Ǯ���CV�R�>B���0���;xIu�����4w�#q�'Rj�nEQ�Q��J�7��{{�$N�����|�2���w�t|�o�v��� J��x�����7o������>?����ۑ&g�i芿Y��5F�=B6��>z��>Q�%^���7�A�]��1��+�oQ�iR�{�cme��7��e<���Q8���=�d��|��S��]UB1��hoB���9b���2&ͽ]����[,�ު����W�c�F+']C�PW�w�(.P)��ZW
^�[�sm��L����~.��DA�E"���=1����)�%v�˪Ԑ��?�&Y��X,�����*�~�g�+�3���e�̔as2�"M%�E)Vm#��BK������r�]�ɷ���[�K��N�\q+<�3��qڽ�:��#V���K��3�J�KQ�~� �_�9�V>����	�IUԪt�
w���%G��G�h�Ad�1}�@�Qjl��5�N�-zj;������š�H5�kq�e�>��j0h}�bs��kw�{*2�3FJH�
k�L�-�8f-��Iq�vq�KL�AF�?��)51�G��?ZU1�G'���.��{�4e	�� �n��"l�ReZL�yѮp���P}�n|�ԙ�7�=�啃��/�˘(͗@��b�����Z��Uf�C�#5�ٹ�ͨ����&x��{�Y��$��+AS��
y�=sH��T%����??��� �m�:��`* d蹈 ��
�4��M�օ��9��)�k��ipM^0�䍇��V� KQ����D�u�B��|8�����=�N�S^ �� t�a�N^�`ѳ���D�[8B��C詮��YX{�8����(��B�޷x�J���m�E+Eh�[[�Z�7�|/���V.]I�*�p���sç� Fz��
�����/e7����*�j���"�ѐ���V��z�d�a�}�^�u�&iQ��k���pGLZ��.z%@Q�<"��`$B9?����>����m�T�խ=Ϲ0o���I^�����N*R$�A�~s�CY��bJ�I:^JK;�h@<S_���#���h@Q\2!e;"�02�4��E�]{Ct�R�PK���_�~N��ք�*(ShTn��VU�cT���{���.!R2�ES`��z;���b���D��܈~�)���@#����Oqh��c#�	��]��~?|�Ϟ�B� H���^�}&����a\�ڒ=����bk�0�:���D�U69vP��@8~e.�X�Dڮn�C/�-���,�4r)�ZIZeE�0H3+�4�'������Vd/^�g����Y��V`���ݎ����U���@m�kZ�7�*I�������UP�_+3���x�c\Cܓ����5�%��y�l�ς�N�N&�$�?I��ӵl��n�c���9G��c?�Mp8���A�1@��vz��U�~NEc�	O  ÿh ��xֿ2�Wu�B&{{!Z��9��/-0�j��xC��O� ���s��̟��Lzn��b�E$J�Z��3���\<$P��Ñ�+c5kZ�*�~���]GOZq�?�YM!�P���ż:�賟��6]~o� ��1��rK�����*�
��L�M��X#>2�_ q���}�U�xU�L�ȴ�rEqw#�֪��N��h��29���UO��j��6���n�_;�x�R�0�-�+�ZD�{H�Ń��1�� ���eⶮ<��-��V�4ځ��R����ld��ɐx�����0W����|r؊//��{֔X�l;|LY�U/k[fs2��I�O1GB����}g�g'��ô5}R�8�����;#�	�y�<b�}&��k}�W���+K���ɕBK��ѠZ$��d�+�Hb������k�f�"7 �����'�0b}����óp�C��������gN�m��S|G$��A#H˝J�&$��M��:op�%�x�(�٨�H�"[�Cܡ%�L� ��yrBn�tχ�lЩ�0��V���b-��2<<Ycz���FZA%B�A��#ٜ�ܡKfk0��VY-�]$�w�I��˯�&A���K'&�Ĩ_92��R@�������u�o;iG�!���)w�3\���d?���^;K�/�.Q���(�F�#^EC�8�|Y��u���F��v86��Twt��*ׄ�����Dw�y)�^�ڳȐoΨ��F&|��W1�#�kG�l��ɾ࿟�7�}Z:�+�O��:[q����k>�L�*R��i#�~�;�~Fm�$-<��j �į9��ڸo�2����#aR���I:_�KJ���L��s�j�8>|��6�7��w�$r��\G�_W�fPMj�	Wo�d$$��E����e����Q�U ��L��7����d��0�w+��U%��ܤ�s [�qώ�x4B�6�k>"%X6�/��FX��>�3J��%�*5N���ȶ����XV��ĉ�T�q|�1���r�9bv�;��f	���hS}����Yh��m��Hm ���z4�p��$��~�=��<KXK���/]������(M8�\���]���=6�d ,bS�/�X���H�cg������	�O����*TD� ��Nŵ�n' ��,[|r�������=0��H�xH5?������r9;r�\�d+!!�����u��� v����|*���ڌ3��DK7��E$���h)��jm�/�_���-�a�^{�t"<BÏ��;YŰ���&A����r_l��X4��������	QR��������4S����<�W�R��G�([�ډaT^ա�(����w{�`v��p�=(7�\j��8}�	F�\	����<�b���%���?���/uw�ѣC Pz������b�� �3.�m�u|���uUv���Ys���<�ݢ�
&��}�,g۔ԧOZ=���U-�f%��j��9OH����,�T	�����_��q��"hi�PQs2��:�}�?���8�����H�N�0���e:3��Ww����_FiVO��؛�S��ד��|��|���G���jo�; o�n��������	����~m/�,�Fk��}[���M�-��^)��p���M(-v�9�-�	ui\�E6YE6�Ik  3���BB��ue��X���c,Let��x��wQ��<�E�c]�#6�U<��p�f��F����c�,�AL��WT M��ÚK䟽^6V�G^f.G�I��X��)��[�_�Od	�#$q�#��V#]#\RFl+���z�eP�`�B�A�� /�5�� �Cf�ڨ�s>��<N�'�ԕ������W�c3��~���v���~�I���)pFCΰ�̷P�OH2����T�?1 ���'��c�e�H�ii�dl���T��b�˛��F��/�TQ��9#���Q�4(��M � 3񔵦�3�����8����@c�}*w�>�_�u۰��lj�ˀ	J�1�Hd��T�g覃Yn��D�q<��
�q\RC[e.����p �8Q����_������:
'�j�7�f����	i�CS��ہO{b�f���n��%����b�s/W�����̕���2ڈEs���y��lʎ�5�"���&�| itB���&��&�Snr�|7�\��l��O/��fɲ��:��mK�@s�6�+C��	���߷?��|C��=2s�+�F�k����X�Yg�Z ����/
��J��^�����蟀��5#�i�Ԯ��&�X�
gU��&X:;�+2������(5e8�X��7ZA�&`���zT���H��5x~I���J�V�G��)x>#:�\��6[�J9`
�/��<��7�U�2̆�hIՅ����gɺeh�����X�=�/��{��$f�sD�@�ul1��C|���o]¥��/�!4�Ex��h��9W�,��]���)?	�����ݔ�.�Á�1Gb�x8��i8�X���ρs��B�gTM]!�� �/b��$��~�dL)0QL���I�{�"��d}���{�B���g�k�w��TI�a3jl�zU�謈98����w��:�N��ڸ��0]ʘ�W����ڎ?+k�=�S�#��R��������6N��j]�*WVN҇6���$���ي�Z׸�d\b�7PAX]n�WbSY;�'���������&���rnH�<���y&�נ&��rA��]�U1��%/I�+���C�ͪXW��{�������k�����Bo�m�����+i��_�+Tu�/>��|�/DKq	�s9l���Ȟ�O텀@Ӣl��K0�^߫�e,՝`�9����F��# �=�����x}Ih �S_�|_x��u�h0�x/�'4]�gW�Iv�ay�����{%d���6�o&�(�њ: i�y�,��Ixd�n�<��s?��!�ן��%D���Ư�1x����ƀ��{63'�/�)L�����;T�l;4|��;r����UXoF�ԍ�x~��m">sB�lJhO�f�^��^�0�/�f9�pW��l�g����7Z	W�R�9�;����E����//[C�Z�Ei���A|i��΢w�����N�����e����VBqv�>�RPej0�	Lbg�ST�}��/t}֊$����0a����#U_����]QXG�/�B��Lo�"�Sf��*�$��4���j��Pu����	�t�\Ӎy�gtD�c5���A;��Ʊ�ykx�����Z3j��l���w�|��c�(n����+���)�Һ#D��5l��,b�����)��F�k.y}+�(���@1��.�,;c3D��wC�p;��N\��h�Sl�`G$���b�G\@�mMB���ixW��G�=*=�J��|�:�A3ФzxvŢ��jшɥ-&�<��簹_x��%�uN4<���H���\&Z��j�����/�|X?	��@��X*�_����XK���n�6&<#�!� O�ƿ��$�*��zrGZ�LMBw��)?���<&�>ʊ��؟���R�|���m�茆~���	t�?��,�3ŷ&F�d�H����3��`}n�$:ql�m�|i�H3������h�~S~�ʋ�y3����b�v�7�<u��o��z!����^�J�5�b�g��pF�c��iȘwYS�h��_'P��V��q���Jf2b���j�\!��δ5 �J�:|��	ؿ�߭	y��ǽ��6χ��4�޻l.8��Z�������H�Ǿ0�Ѭ�Z�C�����4r�Dc|�2�0�~p�Qbݼ�f/��B������`MU��x�� '����~/�bO�mb��pd1���Dx�?�hB Qjs92�����vIY��;�}��(�	fߢx� �Ɓ-/s0�Q����ub�(����b�������J��Z���P)�?����(	��9%"�3y�毆��d̷��rݍ�;Ny��7K��Ě�S*sC�1F�Ai���]8v;���A����A�����P�[ ���_���K� S9a9"�~���LQ?��P�=6�p��t�P����Њ�&29Ks�b�E��x��O�R@�E�uV��G����z��
,C&�J�0@�����pd0N{�g�t�t��\!?��i���M��d���D�I4�q؇
�h?<��eQP�������@�xd��1�t�ް�����:щ�(1�X�Y�)(l=����M̈Q�F=�M�V����!`x*���Y�������c7#z)d1�4
g[�q*������լ`W�����oO�嵥l���ʡLmCʱ-�e�)�~����%���s�J{��Jr
��q7�v||7GӸ���7���΃���)����5B�̥�S���nns>�w[#���T�;z�c:�x7	�/+�6�)�_Qd���[��n1�KLv�Zn6v���m�H �+_��BA�)2������<�}��* �.��OS?9�P�W����a��Y{R�G�K��ºv�b_�{���-B��F2$O�n�t�>�_����A����Kqc�_�y*�3*��۲�r?)�j��C��+�X��MD����܈Ž�y���2b���̑���X��ƾLp|G�����q@F���R��M����*ݑ.A�/o}�*����ܬƝ�����Y�xA!�F�uc�)ЍVk�,�m���p.�Fw��Bk2����{ j:�[J���)*��Df�-�'��%Vv�G�����XA�V$�i���BJ@���WVټ��/���f'�;����x��h��'=��(�Rd��a�7Wpk'��7�FJY� ���p+�9����46;��v�C;���j36��B��/��d�+:7r���Ɵ��������f-�r#��9����*k�s��ݐ(�E7���?hy�f��p>	A�u�$�O�B��#���_��Ew��=�ӛw�qa�(��kt�5���+���5�
�3��5���Qha A�rma'�VS[��L�O�<�6ܽ�|�.��������c��d�=�x+.i���\h,0�޵*�.m7����tƳ�]a�ѿ�m�}���>���{�)�w�if��o�l�K��ڔ7c��LpiT�b���A6Xm�V.�ԁna� ��6L�=v,���H~r�1�П�E�M~������2�Q���|�g��J&y��<��B�J��m^ x���bI��b��WVC]{\
0��=��Yѩ/ġx����H��dܑ���t�����|bY�J}��x	�R���K{*g.DS�t���펝5�'E�s�������J�be�g�Ju�Z&"5��~�r����nб*�S��!k"��FNȵ�:>N�링;��ߥ����g��[M-�ְ��6!�6�L��̝t�T>Jz8p��f�uQ�u�oBe�b���RUL�Ӈ��Z�2�組�dVO{�?�ras݋a��-�����L��?�W0��_O����,i�H�q����ja���MD.�DC�����˷*g��θ�o���s��BQ
�F-,Ѱ��[lv���Y�-�V��;C_
��I@�&��kkzz5Vհ)$�V��	��Y���+�Z��ND����L����X�z���طX��hM�0��1�H�|�m��<��P�� �1��J�Yy�͏��|&����{�:=�ȷ�E(,��9o�aT���6���q�q2>�:��mM��v�=��Gbg64��8��p�-yqĳ�j~�6B��ҏ�`x*z3�*�Y�)U�NBe�I��;/2����t d\���b���B�xs$@�c|�?�������_6b��=Wx�FY� �'�i��(g�bU@�)��?x��k��#V�$^I�l2FK
xA�g~Eaƿ��J���{��}x�aMt��6dB#`�����N#���MRfΥ)�HK*�O&����\ߡ+���zV![������I��`Hк(��	���}�%����8��^�d��`�}�N�$�����g�Ȯ�Z"��+���bκD��M0���J�c�+E��Y�������E+-�`�a�
n¨�K��FP�������.�j6�F��!|�Va^����eo��3�J%DҶF���\��"ML��6�%��e�,���wx���)���%$L�]����R4�!\����G�/ږx�6������8T�{�a��%ڤ��̜0�ȕ,5��}c�ښq2D��(Or����/��HNh�� qJ��d�l&mB�{�	a���?x�jỄ����O��x�!o�III΂���}��2�E�kOT�Q����(�j�Ԏ溲N<�tvy���4_���G�P�n�䤵�B�~��[QV�"Z/#*o8���'�W�x���ޕF, �6���k��c�M���I�OMS=@���}�׽�OF��ws��2�[��%�аFŚ��ǩ�g>'� �����[�E��Ɉ��uo'0(���H��̡�����9#��Mw����1�>�A]�ݖpM�w6u�J��Eڻ C'�ovh�X<���2b5T\�#�[��Ѡ�F=���(� :\��E�n�ʢޠ8w�SY� ���� �z�����C�Y��Y:7��-�=�W�Ow�U�m�Dd�����Ek�"YN~��~+D.Ũh�/'+>��9��{�P}��3m˄�D0����~ѭ��9{�}k`epX�\�c�����w9��k�/T�N
o��I]� �5~8pZ����ZR�/��
��E7Q,���������>>��x�S�w�S0[Ns�KK���������au,��O���n�@�Jx�1�I������!��0�~� �C&JvtH�FJ6��-���V���3��
0��'�Yx��1��~\~h��%*�Q��Kቭ�{)La�YI�R�]�Dͭ��k���K�t� ˁ�F��\�*��g	�[>"u�,�_&��IA�Gf�3
�d��G5���X�}������W�鬆��RGL��<�ːg�5!^�CU�v��{y��K�=��W�dSR��uY�(�'�H�m���@������.�o��������/hG'K�e�x��SS��ś�4{XW"ØѲ_�f�k3�:�����n����9�"z��֙�.r����hX�Z譬��x�Z��o��*��"���^��Y�F��&�E�4,�==,������RJ�^<�<B��#�,OZ��*q2��ͱ�k2T�e���DѦ����UJF��_d�t��SG�:�t��颯��hƠw�w��|LK�P1���R�8Z���H`ss�T(	�C��'{ q0��F\���זWA�2�D�n�͎�@������&�Z+O�F���&��{�[�V��vn�JM�1��Z�8r�����[:�6h���R!�aU� l�t� ��.$����=��92��z��h4)\�����z������%i˃�B�d!g����LgtE���)e����A�=��̉u���RcS=q�H�d~e�y~�y�B4�;���GD�H_��M~�k����>E����"֮���� ��i��C-�Ǘ�zҕ䝲�Wj�R1 8}>L^ Vi�Ȍ��̴��T�d��n�Wv������C0�-��~����z�]Ԏpi��d���eC{����s�h���4�p��e��*����2��tڷ��'�!~ �b��*�1^c�X!�V>ºU�q����V����}�@����h?��F}ѩ�q��A� ����4�2�e3Tk�>��,y���x�_yV�vr;����GՏ�i�+��6R �xt�����85���m��v�8C�cHq�8�A|a��AEJ��e4�+�{�o�oí��q�s`���i7�q&�!�T$�"�{���A_<֡U��|����N��x���6B�L��$�����iy���D&���l��܇�ε�I�S� #�p�$��QbV�:�S4p�+�W��O�9'�3�T4澵��b0�T�J�Z#N,&ߕG�����ȕ��ǿ��i�Z�k�4'��4/G�w��97Fte��4��Xm����9k�x��:�6;�s����9;���.{�_ޱ�=��SZ���ʕ8� ��Mci�T� �X���&NL��(&���EL��K���+@�)��g��0\��*'�M�#?	w�,y_B�h��ݓ�!���n%������2��M����`[�r��S%�.����?��u�3����'}_��_�[��ٝy���@�4Xާ@B���V~�(0�1��c%"ʳ�Xj`�n+�\0�%�Ro�n�[� <C�}m���$lK�M�P��]xV���8�t-�Qz������[�����0��l--W����V�(��u��oo^�H=O�@�-��:�f^]��FJM����1V?��`9?	n����L���g��)l��P.e�`q�I�I4�q����S�M\)H��E�I�X�漢�ї��� >T%is):_ɀ�cE�����&e�J����j���G~�����}���V��5��F�d=���(I�t{@���v*䰰���ʹ�3�6��¿�wq�:ky4s���yL���y�3��/�cka�	F�?��C>����",�se|���Pĵ�dǢ��l�c՜�K8���'\i,�=Z�M���u�دS���E��Ö<���fޤF�c�F+��o���=|��-OB�>w��]���̺����� {������C��c����=��=3�,n�v�\�����M�b���+�۝$>��x��C��"ʻ��u� 󢯯�j�=�JA�&��H��?��P���3=t�8�`h��!�P���Ÿ�cJ}ħJ 0=mD�,�d��$Z">��I��	����Ɓ����$"�b�v�Zޡ�U�����G�A!'g�=�h-`ˡ!�^r��V
W|�ŭ�f�c�&����-?F��
ow�������$ ��
��|��ɗÃ|�Ӱ�	*n��VQ��ucԘ���r���bWD�|G��.�y"\$b%D��E2S�