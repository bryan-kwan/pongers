��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)��<�=�!�R_酎�����U`������g_Å��=����))�m�[1�@���Y�8[��Z�y.����AN���<��C=���I�QKf}�ܨ��
��S�R��;������#����7AqE-K(�{p5�A,!�פ� �
���gX���GIר���{m�Z?��f�Z?�nG���R패�� ��ނ���� �����n�����m��'G	.,�DSoY^�L��J���AP�ێ��c�Y�E-|�p��p���z*�nm��քȊS������`�����AV���J���P�qBt�*�U��^��!eZ#��
l�Z��t�‶,���V��@p{U�W٩�?�� ��Os�c)i�n�!��K���vh�0P�1�}ڏ�n_"q3��:���w|XbB��W ҆�)��k^e�ˎ�Z|��q?��!��-�c�Ք�B+z�Q5Em�����7O�[���ɺ4f���s>�ץS��m)����Н��F?�qm� f4��Q|��uҷL˥m�/ɺ<��y�i;����.��Ԉ�xi�t��v��E6ܖMc<��(:��y��C.��~q$�T�PH^&E@#d�v5��.�u�4^�@�m$P���������H��!)i��^�j�
-�R���k�l��� �#�� -\2�&V��'�@e1�E-+;���8Ih�GP����Bq�s�cϰ(�8�팰t�U(��s	!�!Q�~�v,zc�M�^��i>)���95�WE�(�G?�����3λK�3g���[�����H��`p�:%��Sk��'��p�η������aH��L�Z�6�S@̦Yg�d��Ǿ9�C���B6�����E��}(?w"�ڽ�"�3��b��=���xS(,|��5TSo�fͱh ��jO�J�\��b�]���*�J%�NO�-<k��G�p�P��B�*tW�K����?��}]�"�Bq�R&��
2��u'{cO�Ё��,,['sl��s�(�2Z�i>��^s��7�-x� �7�#��D���uӔ��R�\�f�V�k�}qbD��)��chKK)��qX���rp'�d�i)���S[�KJBA��2��{��ka���;��]���t�؉�0�[cN
���vK��5��4"e �������晲]Ř��d��2�1R#��rF6^_S��B�-S{�i�e�Pf���N.=����o��������� Б/^�oRl�8%��/�h^O;���m���ڝ�aP���w�3��o��<�߄̉��8�ⲫK\髏��)�V�M�=S��N}�6,�H�2��/��YaS��+��:�b�lt�OJh>2�GI���J�QQ�4�.i��'�,�Y��������<Ɉ/���MHw��ס�+	N��-48��,9e�&��`�{��F5��?���O�S# Ío����a�����(����$���	UHA�g��aj�sO�h�:�w
��(i�aC_ep/>^q�f��_bC� �m�i�W=��3����̊J�Bg�[�r�e���c�G��-쎺BR�"wrYN���k�m9�>�	���dN'��N�K_0��Q����|4/���,��׏I�>�r��`6��=�hC��a��S���,O�-E0�����9�I�2(�Q��)g�D6�P2J�"В��f��ԧ��'c�b����7}
��=�V�#��a�"*�Xٯf�E�(��1A��l:��&�nq���]"r,�~�1*�!�U�\�+��q�`�斠��$(SB�v��'�M��<�?k���p��HD£h���s̼>�	���i��뵷t�c���I�
�����`�����F�<M
��+���F!�ύ�X�{��>�2�1����"��l�1���j�
�z�#:�~w�H�f�}�iVZ����O�+��������1�30"L#pc�ѓꦈ�ŐlD|\�,�[�huT�M��c���=�fl�s��
l�g���Z����AIy�^e����A��6)d��ɴG�� *��W��|I$�K����4�!�ݨ1�ζ/�eS�No1�������*�`_y~t�ɶ�Y{������	�a��7bn�=���_�IYT��
�s��m���*��=b'�޼)��`���$&O�?��1��tIcF>7�"�j�"��
G��X��|��'F���l/�0�YV�����5]��M_$SN*A�*;r(;H��S��тj�|�ծ��R�*sf���7g��z��K����f����f�!�Q��*��u4-�lH絎�/�!��{
��Ӊ�E�'��kL1yc+�E�mX�XY%�C�E�	ߕ�](�br ��"�����X�}�f�����A��ݛ�@5Gd̻E|	�v�I揘cL�2\sЮ��r��x�����lAm�!v�&�#q!z�*6m%�
�A�,�M"��2�$�/���X`�rZq������~�M�GpU2E����~�P�}�1��c"A�cx^Z �d	��(ֆA�.��z�Tt��6��T5N=�.�1�	ӫ/���+��+��_@Z&lղ��/�0�:���5�2 �<$���/��㲋������/<Y������-{T�[b�:�	���Y, ������\S���
�Bk<��yx�v�\�	��cUҳ��t���~`؉�/�����ȿ���*d�T<P� #�L3\�vxK��^6�,�4,8������k�z��e}.5t����Z�:�k��i��n�u�ir{����1�;!�%��AL!�����1���1;E��@�#w3�c<H}�<��m��X7W��zOC�|S��57���v�N��� B�5��+0z��(���CZG��\k�8�`O1�HA,ӹ]��¯��UO���U,u�,��O�oeSXI8����Z��zh�=t6��}6�/7��Le�mu�K�������1"��+��ˊH똬o��seBk���=�ώէ��ʢ���Ba}q윝�A�^�c[s����E���@�N�M �~����
��`�c�;@Z��,�����~�u�O@3��V����M[��w��;J�Ģ�����4uk�@��B�2�IR�A����8A{Rx�P�<_�Ї��Wϔ�fqe�%�򼍀���s��A@���'���鱩Ϯ�c��t��m��;����p~r)G�cR��e�+I��J�� ���� f}`�����,���}�F� EԱ�_�A���������l:�s�x��Z���Z�����)�f�ix�b`8�
�_�����b20�<rXr&k�_�>�RN�@��;+�����@Ucg���.[�Gw`]�sA��H d��u \�K������R���z!v�2$Y�9;��q��;�5�<���
�H�N��
���.ɲxK�����-�2�IԒ1Ȥ��c�5P�?�G��(��j��ETkS�ϘۢE\�=cEO�ڰ������	_NJ����]CH����Ѯ�d����$���9p:����L�M�ى(��d��j��=�5ث�����CE���˺�������Y� ]�G#q�J�ߩș,�-������l�x=n�M�������HB�Op$���%��?G�A���N��M�L�/m J��U �2�m'8'Ȟ�����R27��;F`���e4�(�Ҟデy�ź`l��"�(�c[�'[0��Z#�3EOG��A��mNf&:�?����9���pҫ��ӕ��M~��Uf���`=�(�`��W�RH�D����X�0?��<���|*��-��W�H@g��\0S촾�ʸ�Ϯ��&���k�L%k��nӓq}.ﵸ�����h��>q�=Sn�P�Z�O>4�0�%U(�A+?e�2�i�����Ub�s˒�C[�44X�{f�$��!/F/�E����;��펝>������WmmG������~����mb�$h�zϖ�a,٦�vf���, awgڱۢjWgW�0�# Sdy�\	=�sM%�D��FN����}xy8L����/o���1�J��k6|���XC#�:����2z� �{%���C`Ev�ߣ� 	M*E�b�{6)���ӥ�+8���i�I^�	81G$�v���_0"�	0�#�Ia�A�V�:��-��mo�ro06 �M5�!`���FA��Q�v�8��ʓ������vB-\Li�9+����"7F����g�qb�$Y��7=�t��d����iE&�*pF�o�uL� �K�=��}!�R6_qE�M�e�p�8�xF ��eU�N����B@u�6-�)��C�e:�n*�w��n?h��"�9 <z3W�s��n��5{"���� :��P;�Ֆ˽��\�������� �����<Tp8�Mi.E���!�?揮p|%8�e3d�(|�8��o0��GrM��rk����6`nq.FҒ  .�r_�?�b7��B�/l�Ԣ,��e6�#|HT��S}'�Sf#=�ށA���E'�^6�����[�a=�y�i ����~�1f9p�����!K�g����:d��_G:Z.�B@U��6�(�;�'*gTH,^���R[/� A+	�B����iv�P��+�΁ۓ�����6rmwg����7δ$���|_�
<�d�$'�t_��d��V�����C�͛�-�X���_烾5*���N��Q4T~QIv���i�=��Nk���}��i��w�n�?n���5�{=5^��p_*��zc�^�3��̧��Y�Y;��I�����I�<(x5�wk�]
�>�G��+qoJ�5e�v>U�̅f�����_�i��#/a}a��Ci���^��I�KA�A(̒40p_��1�;.�8�G��W!,S�:���u��fs��`�m�A� x����l([��p<�N(<�7��@�D���^�z/���b�F	^B�����&�rѕ;o�>����+_�g����x\*�)P.M���,��F�X`jUZ�\Kx*(s۹�On��R$� 3��H��5ɴ�e}�P��#�o�I�)ؘO�Q*cD�2, ��Yz���Lq-����!��z��T�!�	��Ͳ0J�驽�2�kR�;�m����e�0�X�3Τh $�E�X��^ ���^U��sf�-"��^7fa�y��������)M���3y��#?1^e5lR�ף� ��.I��]h,O�ҘI�A�&E�Dx�EMa�{(U�����S�%�V���/��i��Z�(5m]`I���!��5�;l�B�J�����xO�ܨ ���ghM	rbECk>o�3�O6�Q�&�(VH>Ӑ�+!Ab8_�����o:�O�%�g� ������gf�z�̭'������=��7I��@�FdA�g%��c%��4)���@<|X��cU7��aŤY�΢��G=�K�jP__3�y�@�p���4р���]0Ke��̘��)i�{xo­� �v�R��=ϙ�St`	�I��>�oWM�ʢ�>��%�9+�}n?�l�-���.�q;�1uё:��2+rۅ#���:`���+A��\�u��4|�sy@⚙�ԝ������&�Y��D?ڶA�RM�-����.�I����_���S�)��]�Y��#H��N?��x�����r=o��ԣ�:C��Õύ{�UY-p�C|�8١�+��̀��tk�`{o�BP���f*L��5����E C��-����y�c��8K�Rj����KHU�?�Lb�7*�֪�%t�r�Dԓj�n��f���&BU�hc��U��e�b���Z#|����/E������Y��U�vJ<5�d���pMh�\.�	\������	9�UN��9�S �Z��u���TGG[ܴw��_�����A�c���q4`�MG��h�WI	J�'�U��ń��<D������#�i���*! ,��2�QT�������6!ӌ����vP��e2_해�v>����r��E7��d��U|gx�i�J{�-yo2DuZ��&����6&c����8�����7��Y��~tC{��@����7Z�C�:���P(n�.�je�tR�e�K�U�l8�Bm��ճ�Uxͮ�;PS������H�d%�w�s[��0����N�P�1����?wd��o"��Qc��r�.K?mP���XŶp�,@���=%��Ds��&�|A����d�AP���6�a��eY,C�j ���p���0l`J?<S����vy�����j9h���._��1���$��s$ _�EM)@��(��*�L��U�u�[)�F!�X�w�n�I���ɟ�q�*3?�%�a8
ctkE��l��U�AT`o��-��*�y�ͩ�Q6�_�����g�;�.���D�4���c�H2�+&��)��g�X|�_l��?#f�� �6?��I@����B?�TM�9����:�����*���z�jX�ed�����O:��DѶ�G�
��~N��'��_O.(�n5��1�JJ�WC9T���s��W;�7I�6��vhEGi˹��e�;��]�G��u��a:��-pX2�3��1�.�Ư�_Y����'-#iĮ1���4؏k�%d)L�����R��h�z�	�6�6�Cy@��I�N�����Rld���N���3�$�U���L�y�n(����T؃�2�9�,���f�mK�+zO�&�*��.�ɹ� 	��m�	F����S��������* �ZF�@���@����/��d�ʆ�̡\��G�:���/x�ޗ~&@�����˲�> �JA���x+�����e��Y)����Ωc��:Ȇ�z����d�SX�w�w�E)���R�(�"H�q�3eۈ�cB��%����iP~�ю����&��+�W';��ç
�׬�AsQk�A����ٚ� �L}q顢��-�#����k��7��L]���	RV&Ax����9tg-B"�\�c�ܤ�;���5�Ҏ���Fqc^:��}��)�sV��A7Q:\�r�e\O���^Y���mg�Q��� �V��T	Ԣ�`�2k��ܛv�1��C�k&��r������ْ�E�����Nm�6 �ё���_��᭧p[��٫�K�l�I^[m�{�"�5AV��E�����R�\ஆK�Z3"j��1�f2�/�H�?��U�.J��z����M����r�J?6�u�'&�դ�x���\n�f@~&s֚���[༵�^��B@��ج���@i��f�i�^�����;��Sk͈mg�������F�g��P�4�	�&[���B����ڄW3*�R1��&�^|\]+->
�B	��a#Ӻ9�{%��M^{��^䜿 N.�0%�5.n���}���|�
��܃���;E�9�]��g�@�X[P��Z	���XA�Di�Sr&�3+����&`~@v2��Q�EװU+�ЋY�2W�aJ��-�V�Y�����I5Em��Q�O����ڲ=�Q�צ�Rc�X���$B�3����ω�U!��å�����]���*k(IH+u�M�ę�C���`p@�^slJ
Qz�G�:�΁f�Sڐ߃c�YgԄt�����Y��Eg�3�U���ڈ�����MՉ�d�����rTo�z��A�H�.�0��(���O����O	o�F%{��%����H���4���VF0�w�mb�q�^��O ������	X�aԟz-�jMwg���X�� ��/��U3�g�����zcK�7��U(�֙j�!XAٿ�4�3�5��.�N%^���{v1g̙�<*E!����G�0Hlا���X�f���3�wMz��G�Fa7}׆�kqy���r�2ܴxH����
e�z�S�kiR����Aƚj�Lxϱ)� G�๜MD����8v��\���!5!�@����0Y=�h`[=�ِ��k�u�8�i+M��/̉g�H�[8q5�9�u#^'�_i�Y.�IW�:rg�	��-�P>�V0�-������aH�[��Yӄ�������R��n �p�OW9���9��R闚��؏�WB�c��N:�}u�ow"�R��<Lqq���?/a�MԖ]b"����Rծ�'!���G�������썱[<!G��5�j�r_o��MD��Pe	u���zߞR,�p�#��Ϳ���HM�"��E~�ϋ>{�
���Y��|+r��c��pJl^R����N����B��c��7�l�z���S��duKg�k�y���.���:0��)� sʗM��P�M=K�RJ�ś�2 ���zs#�%=E/Ih�]{L�<�z<�t
���	׬m�4��ó���Я�&7n'<ˤg�|Q����:ٲ��G�kB�z-�;�P,���~���ݫZi�@�t���[P2��EͪK&���v8̃/���^�s�*|�yK�(.F��>̈��H����ntɧ�����ojI*UMhW)�	.Ӿ��x9�7��w��)t�G^���5��8��_��"N�m%q��8����� ؔH{8x���y9���Ԫ	r:X�Y��;�}e�ٔ�����X��r�l��B*Ƴr���]�e�M��z�Z����3�i�ŖB?)ۂ�y/n��J�~wÃ��O$�{�p����?�[���͜�Rw�L^���2\;��y�+S��m��%4~�*t�)�`��h��慁" ���P��(��j��	&��Gh�4Ml3JFEH/`�/)4zP����#����O������ �֊������� k���߆�]u��d�i�%j=t��o H���k;>.;S���6܈h,$�R�L��jq�M����օ-��Hp�3^>����*�&��դ�3��Lpe��n~Yت���K����Fux�^D# �W���|�;�����-U'��Q�@��S��������e5T�Geod�nF��nM&�t����̸n�=Ǿ ��x���2�dp�>��w.�����Jh�:4R� �Ht�WS�[��R�&�Ɇ�~�x��̯0�Vެ�2P�:� ����U�R�[����ma���z��!���bǀ��Y�`a��X��[��ǃG☩����w�fO�:���M	��?'�CHl��& m[p��~�zal#��Y؁\�83��d�dF�V��,���n�9R�:��n���$�s�o�V�1*)F�Z�sl
���;����B��+z�*����e[N��0��P7�$VA6W�C�t���A����-�Xތ�U.\Q|8��n���ln�7E��c/o�N��R���"A�;�����4o������LU��-���9���c�b{!V�y�jG���
�����M�!�1+��s!pۼJT�{6$�̆�N��j��I��&� G�[53��^6�p!�������kޱ�ܔs���2�����y�����٨P�nQ0�Mx�K�����_�)��R�&s��:q�g|�����-�Jy?8y��YR����1��/�%u%�F��N��m}p�$~Q茰��Ge�a����^����a+̌��9�����(�q���/3Dm�[�h�rB*�T�' DB,��Mz�]S�dDN�fu�D�J�V9XRU�^�i)�mH�ͭf;Fŕ����'�`�U�B�~p����l!�k���?
p-P�:�j��ջY7I>7��a���E�}�8`�o����*!�Xh
���7�v뒶���6H(�I��)���'eX����b���=��Au-X��
f������qqB�ƀf�1"�a���p��{	w)J����}{HB$�qU����+v��.��[&0�Ӧ{ud��*e�C�T�X�-�BΪ�62�ȷ���'*y�mQ"���0~�Ѻ|pL#�W%D���K8;O�C$ʙA�	���~#9K���%� B����5j����s�,�{;����߽��
5OyJ@�������Jk���o%�X�5�g���Xu�!_�/}[�c��M	�V-yT@��݂��A�M�i u�D�����e�6]+OE=Ϣ�?�<��yC�2�M��?Q�Hi�A�O��N&hv�c��*Y7\e�螁@694��&�ό�ކ�$Kƽ��?��H��?�@���Р�G'�u�0�~��a�.
_���yn�'=IB`eER�����v�1�.���t�`�,oM9�U�TSV���gB��=�=r�~��Z��|�ɣ�fˡ�����BYC]J>��ݜZ�>�TH���%�6z��|�Bc�����0��D��c��?
�v��J��9ts�JJ�佬���%�.��R�����x.S-�	xs�{0��L>��7�*w
���M��SlR	�E�m � �ɐ+��; �\7��%������ɹ��S���h�<`XucԪ�b���X%>�!<,��]��
=t�*G�Οw�	����gE�^��7u��>~�t��uJΥ�B~�������1�,�a��`^�=�?{|�)gZ�Wp�4�X��=�T7���C�|��!&8�/Wְ �������)�^D����������؂�U����^+ G�
�F�b}f��J�<mf�/*i���Xy����+���l�їݗ��.J�����4e�0�VP�����&֩Ex��#�H,�n
B�<ܲ9Hx����-RX�jl����#<�g����;#Q�]�h� q?���Z���麪�Y�%��+p+l@�_T&$�u���#h��h�2���T ���9�pu���N{s��Ǹ�/4�������kx�|� ��:zF�F�A8w�J�;D�s��Cӣ3`ʔ=isbmf	@��[OlM��D%yR���d�{�sS���"j�t�#���n��$=��l�3T=�J�F�)�9L9��ԝ	�,��M,1v�Cʵ��)-t���Rl�r��~H}=^��ڶ�n�Z�d���-���yu�SH#�R�tP�Jh�KX%/yW|?�]5KN=�q�Z�8zN�:�׍���$	zх���S�p?<'n."KYD{W���6��
�����Zr������a,P�~ߌy�rUP�Α�9!��_-tH��W�$�PޯuH8��O	�{�X�)��{�y1 }��TҦ�ސ�V ��r��toP����3�>���`6
�Â�|8�>�Ln�˨�B�]g΃��*GB����p���2G20
�c��GA��<E6�/o�ߴ�֢��'�T�^�dC�/�^h��A�.<x����'�m��ľZ*S��6E)nĽ/��Rpݺ����t������P�-ќҏ��t�@}�<r��o��wƽS��=�a���g<l&x=X��Vq@,�Wׂ��$h�]��M6/���xc�s�;\��I�r=^���4�e^�iY�KY��lu��飣B�W\�N`�a�sE="�(s;���<L8���,���XU:L�ex1�S��;)&~��׃紞?K��^s��W��^��૗�\SiT��b�����H�y%��,|v����/��<�Vĝ��ܽʹ�3�dcV�\0=氷�h��Xퟤ�݆��sG�b�떬�LE��q����_Eě{�ۅ��U��_�7���%]��_UD5Ϛva`
r/k#'�E=᥯������������R+�c2�]I���&��.��Z$�w�]��8��s��aG��m6Z-u�/��6�d�rP%N	�9 J�A@������n+�Ly�b\�'��3�٦�0㉟q���E�5v�Z"��7���)��i���+0-qg��j' �25g���Ӏi%j�e���W��<vE������@�m!���3���H�bU�0�n�Q*�t(K��^����GU�b�Kұ~޼4��C�j,�����T.���+Y���QV� ̦?
Z�~}�
0:��(�Y����؇2/���X�wu�uAbX̽c��x�M2 c�`,Eio5�9��	�mh�����4����׊f��'C{�(�����sq+�{R��CY��_d�=˿h(.ZS��y�c�?�� ��f�#�vp.�EJJ*�V����&�Vk��ۼ��yҘ�9�{'���"�P7��Z=
<7ZOP�k-�'p�MȻ;����O�U�zS;�_E�i$��4��zf�߸�s�t�B��"�����ѨO���'������.�x�)
ޣO��l��5�5+)��Ć/�Ά�k+x^�"��,(�7�h��%��o�׺W:Q�ޚ���Ʋqd�J����:��g�w�z�k������ ��&AC�����雟��1��p\�'������
�tgu��Bf��Ȑ��G`eL0�t���L�JHR�I��q�����J����;������(��9��l�拜Qf\�Jm�`bK/01Ǡ��n �6��T�����s�E�7/�j��Ņ{��74�����L��k@�Q��|9D�`�YPT<�G����%��������*).��0nB��}�O�A9,z����u�Z��m:վW����Oz�(JI �<F"��óM��l��H���W+��V�4a���Ji��b���g],�I�H��eEtO� (��ޔ
����r��Qֺ�ۊ&J�^]3�̑����#+�e�l�qZ#f�W�h4?��>��Q��XLN���� ��p�?�]�[�?�JFl߼���X�5͞V1[�
�OKH %�s!�l5sU5@GJo�nwq΍�{�����b֓�X@�2��6�g��D(k*��it��</߶�97�%2�4��)uk�Hd��%��k�F��`�$�W��~'��G�f�G���я;��(x"l�|ʷ+�B2 �3�(�I���.O�����a>zj���;�k����:�E��%��|CP���w�['*�)�7�m�fA
�eT���~�њ�gsf�VEQ��E�lRN�5#Yr'��.�@//lpJ��ؗS�(�J�|���2������O�Ƣ9�a��h=�PbHb���������2L"�a�Ȅ�&˔Q>�vp.��mv;M���b��X;S;�AV-��/�ś�S�s��`B�٘XˁA���t��z��ٲl�8,D]���D�����hR?�U�������NI�]q�)�-��.�ynv������x�zj\&?/X��x��D�K��o�=�-�*�Y�ul����ϴ��rĦa���T���q����#�^�;�k#e����E\�F��I���Cc@b���B	SG�w��-�T��=
7���$�Tb���AG3��PL��"�«����`��z����،t���Ql����L �-�t��{)V8�O(`�~,P�k��rեA@�"md�"�j.�1f��T��6�"��[-)��}Y�Xx'lS�Qk�(ð8*��=�u���_#�)��B�������,^8���\�̵��t>�֘,s._��������TB��^W��m!sa�-����_�`ivl0bվT7^e/���(߬IE&�MJ�9iu]1��x#d�R�V��� ��q�m�����2�W��[� �n���Y$��N�P�ħ��"XPz?JW�sW�N�Q��M��]5�.-5鈹���e�c�L�c���<�7Fi�wGc\Q	�eA]��pAb�{�M�T�#u�O�Qz����j�߱p��,���4���ݗ�Ħ��Šg�.�r��腉4�t��VEAh��C�xL��ff�{���UD+��hxc�����}�'����������4*N7�q|�nіw�[:�k�g
����������\N3�p4g�@[��M��s�wi)�w��kW�7{Ґ
���OI|6[��Afo���9d��O �B��]�H�+>��bV��ѭ}h�:
l�R�0�V��$f�<�u/�2
JV}^6��T�'6!�;ɑ��l�a��L=�S��7�y7<7k�ѹ�Sm`�S���!A�B�W8xnN���D��̻��Բ�7�sɋ	3(p2��$&�Cj^��X��G���4������G�Z��� dZ��=z����:W�FZH�V� :�o���V�.S@.�1Z��?�U'+�������Ę7�[$�=iN�F�&țL��ǽ2�������3�7��j���7�jgdaxp<���u�"y�O�^r��5o���\���Fu��N��(x����~l�0�����I���DZ3.��L�۵�j?a@ʔ6A���n۔�!�T�c�u��	�s�0���.��$�'�Ix$F�ʢ���:D`���r��&��9��/������M�Q��XO!�_��o�����8�|WwY�DpSc����>!6�|^�G�փt���2؛�x#!J���:��=��:���1*rh��K��z�g�7s*68���ɘ�_J2e�D�6y!��o۩�].R;���ԯe*����Յڎ��D��J׋.}K�Xl��sK�S}CWL�M����O�ߊ��sg^���h�EC�e�Ђ���G��w1$j�Α�\���^R��$M�����9`��h�)4ne���7���(�ŧ�?bg����f��+.��'��C՞�M��k�?gbC�ljt���!���8�_�̓x�Rpژ���٬�<ׄ��@y#�4+���zHs1�F�V�(��F�)^�Z<u��m��И>��?e���i��Ldg��텄cU����aJS���q'C�x�ߣXt��w�� �Ië��7�����F��<�-�D���
h;��U�4�lw'`�G�>�D���0��b��x��Ό��I�$URo�Д�]�$$�~f��a�wd�+#��K��3ҩ�S�N��hLd ��_�����PB}oA�q��p�]*�]�P8�Eܱ�5@7"�!�q�S�b ,��]��HPIc.��~�]S��
�����6+[����������5'��0ڐ�\�5҉H����}�B�71T�B)��b%�s� \ �̷
��YHθ�2�]�ab�+��џ��@ބ��_�M��AS�$����Yj�I�K�R��5������E�$/���ft�:f�\_����߯�`� &W�!Dq*���EH�t�
��zD�M��Gi�y)�Ygp�]J O�Ѧ����U��6ZW6�;s�� k�Sk�X��=|Z��F�F	�e�>�R�ƺH�C�"3�;7w��h��% ��&�"ƛoG����e_�!��sY�(R#0�j�^ό���!�"D�hۘ��eA�؈?�k��y�b��f��g�A���U"���]��� �� A�>�Y�t2V�O0����1;c`�{S$5�*�$9���T�ٞ����G����Z�ϸ{Ewz4���Q�(YE�éR�0
i�C�>�Ҏ�1����!�V�������,䎣�|���?��!���>�w���V�\�z��,�R,o�$wj�o�����C"F��ف��*�A���d����QC0k4<�K1Q�(=u�/N����i�Åg��=R�~�f$`9��t�����&H�� XFU�Y��ŴS�I�)	<w� w_���u��T��{���q���H�)�Z>�)�?!ա�U�p�vo�����B�K��ƈ׻_��o3��Ѯ���!�m�w��,�d UCFc�1�ė�?f���0��_�����W�����[����б���/N�;@��#�mza2�����A9�3:��֐iAk�J#�]u�����fPt)�&_]�{���VGQ�|�i���l冖7k�F���;���Q�	//�L6�����s�$�Jx\�M|�ӟ��)��m���Qr��\ɇ'��J�S����(s���r.^��O+��r�j�h��CU(��)U�+�	��is��k#�K�莳����$2`_������e�?h��M��{���f�ޟ.�Tn�@h��f��/t�2��F����t��!a��c@�}�4���=r�'��ṝ�Y��:g~i��ۺ�R7�ҝHj���+w��+�{��*�������V=�MU�N�IH>%��h��!�ҥ��MRh7�q��J/��|�8[�X�
�b=��f��o��u��8�n�����Bd�4��&�b��4;\n-?���,��'� V��[=�(F�8���`2�*�S����U��nB�K��ӎ��`������<�r����.ٔ��m���Ȏg������[��l�Ns~X�\�,4����Z�rљ�[��ݙR��j�Cw4��n?�U{UJ}��,�p�@�^Irc{��+�1�"���净������']w���1Y�d���f��׺�L����[��x�Q�\Ny�K\>����a��gjd����2m�8���d)2�W�9�9��R�����D�sD�7<Z���h������YIr? ��܊�"hX�{�SG��84��y���Z�B+HD���N���Y��E�oZ�Qƒ�]��6%	�)4���1�	��rEeᘦ�>��$�3P�H���H����B@��Y�һD7�/8���*m�����C1R��c�g�f�}'��u�6X×H_Ev�S��~e�r�r�S��%���V���x��؄��~�gT�&1,�횪����<�4���x�^��o���"�ZMqhJ)c��^�;�;�3�f���<kJf�� 6)ɟ�B /; �M�f��lHM8�����"��Wd|�?�8#Kn��<=k�n�A����s����,���s��Ɖ6㩂��4���L��
rq-�&�|�?���[��p�n&l,=č�cb��c�o,�D1�Q�8�R��!�Ƭ���{[gzJ�Q�5�wJ�	�L'��h�6�����Ѥ�V���r[`0Ą�M�T#�%��2Y����Vc�Y<~��+4+ƕ6� �ܺ�\^�+I5{�����g���[�X��t����z7�1"� �/g���;��A;����N]����-j|�*[��eS�� nqy��Ͽ�䔺����;�On-iI۟��pȰ�Im�e�8��r�_�]w�h�n�#(QC��茺}��������%X���~K��d$��m�Y��֓=4�PQݪ������I1: �؈�D`�<b��\���Grn%X�ڕ�4FNfz�釓:L`~�������j��Ų���;@����R,�d=��}mY¢т�/�j�9Y
H�G5�E�֔���C%n�
<y ��$V˳�7�)���4=����!��������W:���,�7����J��=�a�B���(o��f�cck��t��b��������=�+��e;��M8�$����Έ�.���O)��CH����^��h�%w~�ъm���O3��q���5����f�_���M��¨��m.E'�I��QRgK&�f���1�OV/��(>��+g��IC�崺iK�{�t��T���'c���-
�b~���z�-[���v�*������[y�䟖f�K���
��a� ͩ0u�n����;N��v0޻���E"�b��;YO�3�֓b��?�cY៊�������z�ol���k2^_LX�Pty�+�� �Sˡw:�vd�����D�>���\lAŐ���V��֝��4M�yAIR���
֭�[b\�]�R�c��,�Я��6^_
�]���W�љ��6 I��J<Q�K��.�#��/n{���ń�oy�!+FuMD-���d^C}���m ���ʫ�<9#�9W�Q��L ���V���cTݏ�o(5��E_�$�Y7�o����}����w�{���x�ؖ�{g��Q���L����»:,A��U�6P�ƒDJ�{+_r��F*z��Ocvq4f�(M�J��KD�F��!����56N��'�\��$H	�,���
��$}Dx��*����E�x[�3���nKz��y`�>��d�"��<m�hF��Ţ*=]3Ȓ�w���ZkU��!���N��K�A����\�-�Ђ����Q�mɊP�*w����N$��EV益W0��:���낗��!n�Ә8:��N1T����c*���FL�[�H�Ŵ��X��r�ds���Y���qB��XD./7�z��F���Hk��\+�<J=���J
���sJ��^����6�m)���}{��'j�a$̽�["$�g��0�Z3�!���I"�J,S�nd���?����@��r�W��D�"�7[�x�Zѱ�N;�;�QY���{�XmQ��7_ d6{������5�U�̵��ѐ����H�i��'8�J���MH����o���f8b8�"Z��G�We}�����q�P6<� z������nx�,E��4�ןCE�PD�1�{D��WI��9�gpf�_4E����!z<?�=o'�[���	���e�����r/V:��dJ4P�ۚ^����bS�ˮ��[��F@��#$�6�Y�E�$�~��j���/���$�����_c��Sy��h��&�]x.��F[�hE��l�*wU\��$��{	�d�#�&�<�j�k&��	+_jr�2V�<OI�`�?d͛���Ц�g��ʿ6��3	�l3�,J�s�( ��5��;�y|�O$VU�w�97����������;�56�D�c���)(����{2n��K􉭵^���<���Y~U �����A���l���݌��:hU^2�%'t��^��m�=��% Ç<��y{dk�3hcZk����(�6p�O6��h��&ޓ�z�y�z��L9��Y��;^�0��#�t"b�j�W��
[3,���Uv�>�<�Oӹ��N����(S�����_�ܺrcZ�6��l���x7:�80�L�`��?���o�Yx�����-��~���w�yNB�]�Z]����..[4��h����!VM)�Lx�E�,@dj(O���8:ܘ�V�a��>�f*����N�^���.��*�[<�O�k`�
n�f<Oo��*E*�s\@���ov	?�@���q?=1	u\�V��B��2�I�PU�5}UX	x=�!�U��A5�h�ۃrF;=hU5��*������,ٝ�R�\��Vbo	.4��49��9��O���عcD`d9��G�=u_��n
�����O�����DW�j��K�Y�29�A��_ �!yVK@������q�j�Dí/��+�U���)����Su��z�kd��;V��-��
v�p���=�,�;��U�ό�d}�@�Z���i��A��" �u��m �Ѭ�q�tX�YI�<hmN��ሜEk4-O ��u��Rbk\蘍������:���� R��n�>�����P&��|��xǪ"�x�f�����ڭg�B�vu6sO��ЅJ/��N�ˤ)�D�P��m_>V̐��]{�V��CL�0o�J�F�V�ˬ����D�#�,^�dG�\&G����>�Wg3�����3\տlӨ(`�3[�FӬX��H&L!��V�D�6��$Z(T?���'���edd�Tґ�?��X��1�_�n�M~��:Ĕ0@��˨O ��i��4�B��:�g�q����G���(��~殎-Lk9,
�/M���n���Pr\��Tt�kׅ�Lz��1W�9�(K7�!y_��p�V�h���>u,�$��u�j��z���E4x[è)k̡I�ގ�P�0ˁDٸ��Z_��>g��n�Q�a�G4 l��>�������*쑴~��L��dy&6.`c�EY0�O�����6_�ʉ¹�O�C�Y��~b�0��n&����fb�_�W�`�E�zq�3;��-��1�Y���Tي7,
���nX"]Q���a��81��ߺ\l��=<=����aS�)мxt�����s�4��EM#�+��`kQTF0�Jm�hD�Bd�'�x�\.ٌi%E���S0R0�^�uga���`�p�<�<��	FW�حgPK&w��0��0���d!Цܜ���O�@{�N�0c{�r��7L~K���n�Hn�= >���|.����Z�+�j���E�1Dk����Z-�+�u����"�� 3���6��ur��Yɳ�g}ĝ�a��d敏zmS�fa̱Ȯd��7�J:�MH��X�a����?��*06>�|��J���	�*�%!F�76Siǧ0^�Ԋ.��C'iέ�3�Bj�S���Ѣ�ևڰ�}�5���>�R�� -�g����\|B5����e$����ʘq8�:?KP��I��L�ʖ��)@���`ǬI%�vV�5�]���7�(����o��ߩ�_|Gu�����l�/�6�J�O�lQ������� Q�)�g2KOY�����7=���@�P'f��ۭ�R
t�8����M���n�e[���R���������c�'p��S�����n��)�T|�f�oe�鷢��%��4�`�+�+n��l�9�!�Cb���)�2��t.�H;VI���Fݟ�U���HK� =!�W}2��={q���/'�v�e;U��
 I�J�V�d𑎆�M�_N���j����zw��B�hh>��1���by-��h�m�gk#�$=�L�Hi�f%�����0��-1����a����1��*(h���A�����,ٸo�4�t\9�?�5�r�A�~::i�rM��y����sؙ̼��bN��<��5T�	F-H�o�Z��ĻE$��)|��]���'VL���TcG��S�.���k��:k�O�$�H�㯇S��l����0�ڐl*ᘞi�l�1���+�^?�H���X�ǀ��:6���B$�/�mr�B�d#�'��P���M�=�g��dL��� �ݾ�:>�E�z|b�Ic��cwL~��#�{u�y�6��y�Zx�m=�Bx@�����A�S��W�to��S�X\����`tl5C�5N�[�f�Ȕ�5#��@N�ͨ��@��?=w��Q�&(-�-�$��.��ƴ:��lˊ.�Pk1�qW�!] S���ig�J�i	�>��	��JKa�G޵Sߖay��:'}���R9桠,�r����	�4���A��9�c�V���' ����R�2Pf�ˑ����B2P�0c�L���>�#�"<H��skt�{�1���ݶyV�^]s�F��'O��Ӝ�*|K*V��}$>��ư���y���rZ7����m?�[p�~3%5H�Ʌ%$�I-��z��	;8w|�Y\U#�3ӥ:<i �P���l9K�튛��sBI�ЅC�d�8n�X���cK������M!vY��ly��2��M�ܰ_Gv�L��C������p���������RŜ!/aÐ�v�U���D�(R�^�̈E�Mn��Xݢ�6��56S���ZT^�׊��8��+ʢ�<�ǿ��M�5�����My��m�}��'Ms%r����q�U��t�߻�睇'�(#aS���j�nraB�k4[��k����p+.��nt�J��ڀ��5��E?J��m�av�����T.��1�ɫӡ�>M��}��0��oR�����oس�&eIRoVHZv�����3[s���]?�c��69�A�2���b���[��?9(ڸ\�l8d���(����c��?fTy{4��y|<��u��W�'���g���+/�m֙'�DV�s|	�`{����})�SG@����Z��BBA��'��r��D��M~�3�{�R�>[cy��J(�]�t���?VPw��5���Ð��F ���9u��7�#S��vL��e&5�kzlWT�^��`h����,V�&��<����i޾�n'9}�sh��YB�+���v��].K������B02�3,Ư%$pӐ�ƛ�;X�T��������[A�Dh��n�����'�Vv�X^��.�N�\K�~"/
�+)�\�M�$R?�X���B�vpq�C_OZ��kO��V)YV�̖�D�����t���S6:�PSS�=yP�hdzS�l:=�$Ƴ�>A���9цY���d�Z`Hq��6�eEhc�}Б�_�![H6b%�_�.��z��rS�X�d�hY�G0�Z�>�+[��G�i[@E��5��;G������|(oʋY��F�E���e�0�����:����� Eϱ����B=W����A�cb�%X1]DD=�s�ms�׊6�}8bÄ�<A,�(�F�P�!�;��A�x�͝ 4�r��h��K~X�\ko������ �/�賯X���>S�����-�eh���5�ް,��Ȭ$%��}�.���lQB��}Wi.����ִ�#?X@3G�>y*(��m�偤�H����3���'o�.�z�U����޳%��Q���� �l�#�A����ޛ�zΠ��wxϚ�:������Pb�LAi�aU��� .�vD���V�X,�� <��}OR�d\�8b�����8�\��<^�������;���;Vsy7b�JC�U��~!`��!���ˠ�:"@���c�-@JZ�i�/���)��W��#T�B�[�̺[ڨp.'U
�F[� >'�2�\�l�����bG�P�ߠy�;^|~!z�f��m�� 7i�K���5�_��	H4�bt�]?��U���"p袏/�1*�A
c��P��BU�ƶs�����������\~���L�de�V0��r����jQ��0g'������V�,���9+�e�᪅5IiCWԥ�4ҭ�X�av���8W���<�(6���!0o��T�^�����͚g(Jy���"�*eN�+:�=.����Q������l$�}� �ۙYЍJ��'\^��e��z�:�3o��¥%E�oe4 ��;݅Lg�"�Pw���Ii��OջW��V�ҷ�D���*��~QA�}&5r�D}�sE"*@���Oڪ@l<]8E_R()�篧BZƖ�ć}@̗ؔ�[y�*|]��_�nP�I�1�Q kn�yГ��L_j�����Hr�w|�1O�$dRI���	=�QA\��&�b6�.�U�Ul$��rc��>�>�ž���&tk�!�`�&����!�S,Y��[��3�MCVr���E���N/�95�O�8���)-0�Ez3�*PQ#�3�v����J�O���d>��r�:b�<5`u �v����1��0)���r��X�����U� r�N�l��%&m����Z�~�O<�]{�s�K8���=�5:��s:/� (��brm��7���h�Cے���vb��GJB�u��
�At�P]�����`j��%Tla��$��t��(�1O�]��>�[t�^a	5�����T��C�nh��B�bI����� �o�:�03ߝ�,��bE��어uHs'��+p�"��vJ�_�&�h%)�켋��mw���#��:�Z�o�R��fto9�3V�����+�l�uY�����I=�6$�Mk���<�u��%B�`$��˴1�~��+�4�DtW��s��������%1.�+�-��+*�p[&��)�In��Ǝ�t�g�1��)@�1���c�-HA`��1�8���/��-�]���#|��c�
*4'�s�����f�y`�G��(2�4y���ƕ?��7������t�a���:K�{E�R5�|��3��BZ���trL�cl�RxR�R���4g\��i^Mn��:�W������z�`�zI�+��o�0e�������P���`�g؏���]�rȵ z�p���[��!�H>/� ϕYl�*��C��-Goq�ׂuHC$��W��b�y��x�2�7���
uO�F,D�(K�Q��Ɩg?�{�����]w䜝�|?�~kW��^��~��
��8�,��!Y����=��EK&%��Ie����~�oǋϜr�M��L��:�VL܎�+���%��
#�H���.2�m��6W��.F��熗��Rx)���_�Nb�҄N��`��K���`T��_]�<�l9�]�J��y�f�_�a5�R�~>��?wR�!�^7�\Oc*�' �
�갆�J��"kh8lA:�iO��I�y��@�i �0DB#�Ϛ���D��pk.��V��ڢ�Rg��̤�>����ȑ�2��zY>��mXv?��/f�jzn��*>�I`O^�}`�(����7����|) ��CEP��Cn���\��PN��m�T�qcu�,]�6�2�A3d!w�X�����k��1�䱭p�|�6�L^��3�MԯhK���b��w��E�B��V�M����i��"ZT��>�����m���Ќ ��}�~N_����A�������,jA����e�Bw�cM�_��
ϼ�v�?���a�} �6�jL���@�{ղ�K�vh�浞�?�c:��Q�*hB'��t�
��,�����Y'��-�Mڄ����GJ��~���8}� X�Ou\���^L:o��ͻ��/�z��$�;� ���&I�_���8��3��Ӵ���QB��6�����l�F���Y������:��:�-�O��߈t�������)K��(��8v/��������-�,N��Д@�3�.��A��e����f�E�-�f�O}Ծuz� "�]J��~�潉��2�s��4�~u��H�t�)%,ZS��%�����f��$<���k�6O�y2�Y��bB�'�V���m~�.˕�];R¼�QJ/�U���vO����l�>��� 6�1����Cѯ�	Ξj��i����f'�T��V��9���)�֐�?� �)\A9��=(?��K�x�\y$�:�C9��$|�U��KU�ý|�\ ߿΅�+�
fi1���lPP%����[��眈\LB|���q7�BG�W����ґ�'���G/I�+Z��HRNu9d�r��<����L�[�uL�{}'�8r�Rs�̶���H�Ҳ�-����ۨ��p��Kҙ|:w_ngm�$��<����«��;����rHs�wS�=�ߦ���4��C4�xwX��C�+'@v�l���ZP��"�����,����(�xF#?��vLM�Ot�Y����v|�KBN;^��DJ%���s�O�?4z��k�#�7t�V@�7{B�_�ț0��g��0� YÕ�, !��r��t5���Yw� �=Ť�i�����=m�Øpw���!��a �~��F=��U ��@�k�E�k@]@L�s/70^@}����[� �r��rZ5�J5U�<��>
���}�I��;�
k'�i�[B�N��\�너TAP��fhB�ţhI��6yR" ����嗶�VQ��&8��!Q(fh� ���r�����x�Y�Y�ɒ�F����(��q�����j9�G���m���xs���2%�^�5$j�H!%K�H�3��	�P3�6v'���Q;5�%r�I%q��d`��O�w:BD�Ǿ�In�PuH��8������+m<�g��\3|���8���ԗ�*�J�'�9�~(?��N���ۇ��Dt�\D��>� ���Ϫ��]*��e�*����Wb�!dY��Yh�6'�(d"U�_	+[
7�ɟCH��0�u˳���O�/:H	���6Z�Χq�nOZ#m&ސ\��Q���׾�S5�uG��-R(q����+�q���K�(�ߔ�>Vu�̰�^a���J��=R�nF�o���hs�Fv5D��Mx]���U�Mb�bGʵ?<��-)��x�~|څ �.8�Q�,�vOM.�haZ�(	I}