��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����{hi��7	G�����|��4/���YEs��Q��H�9e���ϒ��(��t�.�?�ѩ<�Փ�<�Evj���T�����B�ݰ7� ػ�3��p�����D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�������+�%ix��;��-���y��6XM�F���
]8.�"y5��[S��I~o03�v�4�W�����x���W��>!�3�i�/�T���Q\�^u���?��bUr�?���(˒������#���h������rF�:�8];A�d��Ӻ�X�{'�� �%�]���������N����ě���������ҍ0��^�K���lʁ'vr��/F��7S
1�y�P�V����,��^��:R������Z�V����Y"��v�����Mv����/����1��9r�} ����N�r�'�E��d��l�+eF�V�Ɨ�(��3�=u�c��@Oe+|�U�ve�̈́&3��Z������I����^4�o�B�'ì�n��i�{uG&�cN]�v7�B����K#�9� �qϏ��ފ��U�Ok�x��4��G�e?@��KI8�\+;������@���6xr³�ѽ�$L��&��m!���h'�>q��qU�L���2��N�-^�?�{���z�a3��3F�V�旹t���!�湢X7�z��Y̐��1���v3���]I��x�dV����K:䢞S`:�I��0u��Á��)��?��'����]*�����[�VJ,�v���%��v�k0���A�3+�I�3{�p�T׳#Mz���	���ת��Y��\����l�Vq�'�1�N[g���hw1�)��\EңE�;Fr���'�1V��ѓ�?xI�@҄v59�²}޻x �U�W���j�o��W;�6���pS�|�?io�f«>��4��c5ev��U�Ȇ��)�sqfX]��;�����rL�6�%Oܥ����oL$�`R��\.f�n�$ޢu٭	B���"�Z��]l���~
��>q� ��k��4E�8v+9.�pD�)#�dq�I0 �V�0�����S�t��-��үj�Y	���j�&pR�)�j�
��;�&
�.>_L]_aʰ���4��*TΕa���Ζ҇w��� �%�W^}�)�ABtG��d�~3n\�ؚT�J��)3�����,(��.� �ٵL��N�'���AoJ,�RΪ���푧e�o<�ɳ��	5�n�wEG$`�pD�Z+���N@�jxr'ݫx�_����0R#��ѐ��4v���W�4IB�����x��[�IX��27��U�:������(���C�,J.o6�d��e:�A�PH��K���5�c°�|0��~	�/�N�S��X�U�����䥫�Ҽ��x,��Ӑc�@���q���rK���a&�Өj%_�1V�u\�B���v=��F#ya��ޝny�3�C���	��Z�E�?
r/x��p��ob�����@vq1�Z���}9���G��TS-��'#���n�B�Q�W�[�E��������m�-�v��v�.>�I��Su�J��˾�m1��ц1"��	��g���j����o%<����=v�	0D�SE�&��%h1bl&��Q�H�C�J���� nġ�%�X���3�Gxz��&�i��l��-o���isl-��VFB��"4`��b�����B*
��^n"d�G%#X��?��l���J�%�K�Ə�<����A�,��F;��`ȅ"$��)Ƚ��bamQ���\�����Q $�L��v��u�XT�~ڴ��3b��B�X��|Ĳ�����9�
�Ɔ������+�"03�.��c�����2��H$B3�q"X�����՛��U��O���My�w��EtR�xW���+G��"�]�YIQ��,w%E�)3�ud�d�\�'Q\ɠ8%�!A��č���[�����H���9�i�H�:h���a�ޛ [c�3o��<Q2+��T���]ArL�b�u�xG����"$�M�Z�(y�q���ƾ~�&��A�bJ��g)�kF�c[΃���O)g#��~����q�h�!{��˱�vb���}A���I��^���X���5���6���vˊ����5�	��l`�A]���)m"A e����0���[�e.���nm��4_�'!�Ш��\��N��VJu��x�11R��n��H~�۴9;-��80�o	Qj
��c����lD
���*��VT�z�P�"tj�A�,?$�XĪ^��g��S����[Y��/�1N��.]b!/��k���,
6y�#f��]U��D���Sv��͇��dL��9 ̛F�]_�ݣ�P_8郔R9)�;��]E_<��L��1��Ҩ�px�L0$���Zv�u yU�&F�0+#�����8��'Q:�<7�M{�O��)K��=���>����F1ͭȱrY�)�q�]�dݍ�>%����#�n>�����#�y#���|��v'ri&� 9��LG.�;��Y��p���c����D����_ɼ�;��P:A[�X�
���mP��U�]��>�Q��t+&`���ۖP��!����W��3tF�b��SW�Svm�SK������|�O��@�1G[��uB6e����m�u=�P���%�Z ��`�>r*/$����!-4]g�J���_�F`�rᏄ���#�����j���r��q�˼Xj���<HU��Il/�`�P΁���E��Y�H������<��w�|�u��G,a�݊1<�Ou���f�O�m��Nlk���/��A������#�ww����3��׮�I�NR�n:��Rebk���
[/��P��'�>>36"��+�~P��7~����wl�f5?�Sk����Vن���u��D! ��#����!�������&����A���Ȭ����Xr߼7�.���J[I<�N+W��痺A���:b.`��Z��W�_�%d���M��A����{?y�p{�l���9A��Ù<�-���w�~�0ۖ��Y��K[!+�l�}�_}<~�������hc�|�� �vn�:��=d�f`8܇�ob&��<�efx8ڀLUf�,�qq�e#E��jw���z-���x1��q�7w�ܜ�˱uv��&�J�+pT�@,�f��bT�oz��4̗G6�������鷑L�W��e]�{"9nM��O2
f���CB�С�P�
yg�!lYJz�u����+�#������o�H�i�Tx���%��t�����x�K�MC�xa�Y�f�	!f�^n��M�I��f~%f@sh�(�ϯ<�T�WP- j�/�Q{���O��OIu"�-��������m���ݱVx�~��؂�3d��W.���"�Iy��s��kT�Jږi�6bl�\rl;Jp�cΣQ�+*$�)��w�q��8VL�{�,�}�t��g�;[��m� Qj{?e�s�qѓ�H���f�T�]0���k��O
썺�Dp~��2�3��2=��A:�ۛ�p�j����4G��/}�����LX�xe�Xo0���u�4��m)�=�6P�߷�E@�H$z5��ȝ��qSG��0��G�e�%}S�c��\�%�.�[-�o�,���H�1�h�di+���Wn-��z�'��cˀ�Rb~{�m����G��D�`��C(�Y�����g`���ڢ����-�q �|�ֹ���t���(2T�;��P�=1�E��"���h
ŵ���ҫEM�:�A�TOc
��m2Ek:N��U"H�'���I�M�jb��P�B���	�X�� �H�d6Pk�ɧK$�Â�905$Mo������0{äD�ҫ�B��$;�(�G�R��H�y˰�����sЉ��}�� ����λ�t�'�-�D���Tk�0�Y�x"�ޗޤI�pʄ���r��d�6�m�ϼV���meA��6��$��)���Ka�=�
M���Z_�=k���	%Oi�v�
��>��T޵M��T31�R$z�8��|m��b�5�q�4q��pqVG�\�\�]-���*An�Ш1B7��z�u1��{z�&0���ya>�}pfb!C3��w�����vP�چ�yꝯw�{��x((¥U��L���>�r�}�tU�|8����	N�� !�o_W��<?���"�������껭iZe`�m?t���.g��-:�~m~à�D~ض�)|����H��'�ќ��>S[+����96��(���%��Y���5��&:%)��4V�H����I������;�����-6�%3abSm^8������o��T�nё��2M��siB�2j�۶ԝ�GG��C8��׶�'�k�	2���1.L���p�qRpQ���b%���)朐���D����������P^ђ3��h1����K���}���-��-�_з��l	�J�ĕ� �8�(�	s%0NrI���X	1���~)I��.ռ^�7�H��E:��EoTF�`9L:�&�ԓ�/�q����?��ք�YN/��Ph�9�����l��UE�:���"��廠PlU��Z���N�R'�d�����[���\*j�Y7�')���f+S����U�q4\^��"B�����|�����<��[��kF�*Y��s�U:N3S��@���oM�N%� �E�� iЌ�����}���WHufs�C�T+�`N�ʈ%�י���:���.l�lK���.#r��7wF������1�P��*{O����-�훏T/���` ��qK��� ��_:Z/{���4��E��i��z�'��bS�h��7ƯvEN'��&BR%�W�9�~�pm�v�ی��x@��"|�J�1��#vǗ�cd����
�Q�ɢH�ʆ�7����d�����\r�A�L�smc�,��w���N�2���U�Z����LI+ �D�|�-�^t�%zY�~M��bI���q�=[R�A9���PM<�9���P�m^�(���(�Z��ڪ��C)�hj������:�f0Os���R�z���Q7H�_��`Do�r���"�#���d���v��5x�hHo�3�U*��A+�|X�1��� �v0��X�é�i�2�1�j_Cti){��1f��y�l�r��v�KaX�iV-���Ƈ��LxlD�ɽ(�*�yХW�4DAܘ�4>2����n�(��+����(-c��L�T���a¸U^-���� ��G@c0]��+��ۑv��1~��M�h/�4������b��KDm�Z{{�Զ��-e^����}b����D�s�Rg��*0уN��J�_������
0�/	����X�p7�����N+�
5x�]p-Z����'̢�ҋ6�����kue;���H9���uC6�A:7f��+�`����"P����Ӛ�e; @�E��9w�t�L�	EЪ��⑈Z�n%�W^[�4�����EU��M�0����`YXb�4D|8ӊ�T�޷~)���|{�l�G�p3��3���J�Z�����埑��w�|��(�'B���j�|/g~h[p��!U7z������EtmT��	�%'��_��z^<�z�e�Z�?��qTI����B����c�{T7t��|��!u J�l(S�,y�xx���'b�Y-�#<Ѳ''�f��Z�dAZh�%~pz��&N�踠fvF���#O?	}�?�}�	�3�W�e��f;Q�ϥ;Ш2V��1"&K�u�Y�_(�������Y��s
��y��,����u260"/H.�n}����ږ>YZv[6��j�cS�����:�K:W���M"j/HeH����ǧ�7x�`]��tP�ذ	p�~��ۦ�����oւ&���<���yc��}df�^��6��4̏�i��(��l�f�@;�Uw���R�3t�Mf��9��u�6����]���9q�JT'�v_�
B�ص����Zt��Cc����[,;�̦=��`�3�CR�B�b���5!�ܦ �Q�}xI*E��Re�~�5Dxz��{�$z ��[����th�x�m�uܯ*��/P$�d��ކ4��ҷt��r~��n¡�@cK&��,Pu)�b�y*4�}2ڲ���_d,�C�&F�T��5�֯2g�ۃG���cD��m��X4d�dE�����[�~�/��q2��(0�;M�z�h�D�͚�ǖ�Ⱦ������{��sگd���i�)N#������Ģ�^M{�����r����il�����$���hX)��\� �>�џ���٢��sp�U\	��PY6U�4�li�#)��.��~w����C�2����(�w+��蟣��Bi�Tt�'a$�N���I��i�4��-��љ��!���62"xS8�"	j\;Y�=��Rn�4����=�1�86*�Y�VX��V�9�io$E�Oy"�K��
1w�WF�J��n���4H�wAY85V��ڨ#�U��'n��7��y��TW^��cx����[�D\�<��Y.Q��J�R�lk�WX��?(���h���H1 @�%OCFEͼ87�%nM�k�i6W;�1�E�e^���w�0�������r}뢷���k��q��N)���Ɇ�1���:ZgX���
Y^(ɔ6K?Hp�_��wi�3W�S�L�6rp�W��v���D3\��Zg,���̼A��M���͑�f�����1Ko��-$��U�����~rH�Mڲr��B������D�'�O&�]ڮ����wPD��������d7|�[�W������
�fd�*@Zd��.��¿�,�@���`΃E��A,� �[Κ����Ϳ��#@����*e�X�����-/0�m���Sj�����Y܀2��^޾y��1�k�3�u�I�tp�L��I�G k���;K8ۼ�8���Ͳ�iG�\?��a��w/b}��Z�j�,��wX+dΡ�8�2t��E���\+��K�E=��o�Į��(C����֮�򘛎!�
��_x�W�>���;�&]�X�MWV�Sm!֓��M�F}q�yQŊ[G�3
�mY����A�����u�Em��J���5�us��>���и��~��3c�x2l;΀28���ȇ�q�9�sE����^��qF�^殤b�U#��7=��l��J�q�#I�}eD�����uK��O8L�B#��R���Wc����m��V��4�>��?��Ļ��} U�� /��,�_�2��/�-F4�����Ke���b�75U�Xe"�F.0�V����Eo6 ��S+�Z~�B�3��z����﮷�g����8�ܞx�>d����|T�߾�6���.^bV�o��r�+b�K�؛v!9
������w3w��+~�쐃>��7�*�P�#��:���ǔ�I3]��N������u��?�Ǡ�T��0t����o7�l��'������*u*�!BW��?��
L9=/yw��%ڛ�0�p�K�mFl-���z�|D.��آO�����+K�Gq	h�;lj�#���pN�W�s�h�Qq7��y�H��y�`�[׵|xݽ���P{�Y�4D������(��=��P����KA��璓��E���"�Lb�u�����HM�,���u� ,p[��p������om�J��a�D�`�B�؏>Q�� ��(x��b\7��Ѐ�i3��YX���ی"b�� i��5f[�y��kl�?��nGkf/Jl��d2��ĉ��HD�.��*SWET/���X�K��
�AF����	�A��5����:�j�iI��<�+�MU�;���uyҐ��;���Ƙ���&�+��)�����)A�y��RBR��u�o����Ke������4t�R�T]���r꒳X�6�	sȓ�jP�W�}�}���NZ�����C���Q�g���Ձ�^-B��D�B�)�=,D�ݨ=O�����l1BD�ȗ��5�	6� �l5lĂɲR�<���H$��N�'� [~��:�'��]��n�}��p�����paIG`S�Y�>�4�`��j<ܻ�m#HD.<��S������3�n���T�Y���q�Ά�c�d|��d�=c�Ton��}�W���y��XC��9�U�;\2��������`C���H�N����q��Ou�jC~D���c�1Il*�X�	Z�����G��YcxL;���$qa՗�-�.9v���	���j�E���3�K|� %
A��b��$j���J/���cv�c[Y�TfB ӳ|}����>Z�CSN�� ))�03����9J$��@�O����!/^�^���7B��?tіDL%�P�Z�Ob?Lٳ�3��I��n�n���	-�BL��@FgM�[���|6�ӵ'P�f;�"� ��E�g�,2q��ڰ6BA?�R;�4.x�Y���l$�U9���e�orRV��M{��}���U���rA�cm��%��!��V�����AnU��P�{�*��Y��~9Gt �c�9�^��[�k���U�U5��em��x}�˭
�LS�@f�$"ʛ^�����Q;ۋ�����R�\� ;�87��_ώ���`��z���Ѡq�!j�C޹-]�2$��x ���tث�9���i����0�j��X%p>[��������W�%מ��v���[� _��(]{F�L�_'����&\�����.�[-���5�`�Z"���/�=/+Ln�8�o
�����G�����=kۻt�%���R|�ҁ�j[�3r�߽E�<fǇXu�̼R�����/%'�Q)w}gi�kdC&a���d<�Sd��,p'�����"����A�D��&a{��N��_�i!�b�їS��R�tIg*i����W��ޗ0��~�i�!b'�[Gb�����v�zR�{� p 3ۻ�����ޣ>�L���7<���ρ�T*� ��/PDuݎd� �����-v�T��tħ>�i��Y��t~�?�jE@J�zm��3�B��"t2��&���-���]ן�"�!�߼^����Wvܤ�AL�EQ����a��b|��$�,0	�c�pH�OMS.�)���6p�-P�D�g��`��`���*_�@��{���t��p��]�4o�\
���VH�"�դ�ͺ���Z����e,,����m�ǆ~Ȣȭď�%��&/�� 7�їN���������!�@��&yd��~�"��:��L��V@)�R�$��s>(�R�
6�m<Z|��c����&����'�0���q�|�4eF�c����`��l��p�P�F���J��8Ӯ(3i�/ʔj�#Ba�v���Z?�easLH=�Rӕ	��r��u!�������\��r��h�i�,�̶��S6A>yͣ�T��
����mm�Z|�4�y�������,�lf���Ks")��_I��5u[!�;4�^�'b)� ���1l�}�,AO�W�p/tuq։p���Lb��ޅ�<6/�{XK�^f�R��P=�|���x?=6�6��WW���b�Y��K�`�B�Y x)=��ؓ�3
���6��n�&q�G��>�@�7v|'xTo[�/�ݠ��E^P�&���2�FǮ�7����J?ߦ�4���ߗ쁗���ER�ˁ�_V*�ȆP�,ṕAZ�|���I��/v�2�T���E���`C6`�\�����zy����}������*�N�,L���K��I���&zśb�����;Q&%ӭ׏��������&9 �vd�&
V���"ҕ���g�+&d����|�����mU��o(����=9����pY�9�6y���Bl<��9	�~��c5�x�q�+䎹�(��0�.�od#c���;�'8����n����W[��?�J��"8m�gVE����zt{�5SӝeYo�3���ps��
���D�zS0i��sSg��>����/ }7�K��T�ݕ�P9���:�$%��4Z:��&�E
eO��<���o������NO��)r'(� >�Ή�|:4C�	���`z��̍U���F?��2W�SBm΄I��J�����_���p�񟿡x��J��(��f`�ҵ��	A>!�y��Ôu8�$N�p�t>�(H��X��i����c2q@r���պ���)��.&p�-�ϥ/8+Xv9�K/2V�����$6��m�^^�����p#�˖�u�i+�� #�hf�ah�Zd��5^�����^U�����z�~Ε���XZl��^���UR���~���{�8�k\k��8~=߷��ac`��;�������`h�������T ���n���_�I��?>BR�`���kŹ����~��`_� ��l9Wóu�j̈j���d!��z؎r�짨��o^V�|�pZ�& ���O�I�!FkH@��F[�2�{��bjFU4�Y��Os�@\�f�]W%G��[��]�WHb�	���Es�y-���
:8��o	� *�ZcP*�Q��vy��V:���t@v�C���q�SO�2�~Jp�\ �����E��ֆ�㏔OQv8i�vY��4A�b�P�0��t? X�9h��Չh�}�	ό]g�C�q*{���x6*q=%�5~��i�����^v�/�Z�鬰c��Ȱ�(��q��n<���t�^�8r|2�W��ш�A=~b�K���P&� �X('\�%���PO�f�Ŀ�Z�*T=V�}�Z��_��߬�j��o|n�tK�T^-��˗]�O�:8��{k�l�xZ�[<Ħe<���K!�FO��8N�b��?��������[��{;�)���A_. �}�ڀ��΅aO��>���F��ʦ͍I� ��%I�]����c��R�������/b$;���e>A*�\|_՘쵪I+-o�����d �GFk�oi���Y�8�<��T7Ͽ��h�	`�`E#��p�9����/���v���rb�F!���?D��ω`�
-
�����N����=����1W(�J=)|�n�8�>wks��Q����0�WZ�B�$x��:�dh�*��Io�f����Be��#!��[V_��\n�+���f� ��Q�{����y֩o\C�!oG�)c+��1���ח΂�K�)}��B�з��R��łщ+R�f9�T�c�i��j���Yqۧa�[�SN1(|�|0�Fʫ좻<�P#�i�[�����WF:�L�k:��ܥ��v~��Fb	Ac®��F���,ҹs��{r5me$D9�I��Ț�g񺦾cPyӱ�?����z����`�����x�P�����H-~�P�?�7ti��^vx�*h&ف�F��Ŏ��}#f��N=`�עe�U�]��t�ͯC������ū��Y���N� Ck����� �'42����g����|3-��}�-��6�W�8���ϬA��1{�
@��ŪeU��H��Mr��(*���8�S�J!�8�!*�W/�X�rXq���{%	��#��J+iնN�1�jg�T�0���mA}_���Ӈ��=^�!�s]��ڌ$�_6o�4�x�=JEY,7�3�e:F��Yf2�nX��T�P(����,|=#�n �w�Ck��� �>������A�S
�~��!xKX���6Ν>z��Qh����AC�N�{ӥg�^A�I"��ܞi�Ff���b����^7�-�L+K��R�֠�F��wO}N�����9*�BRv3���j�.$Q��G�6̇E�x�h�,�d޾.ɑ��9�����t8�7��lu�5�}I}jdTj�+��U�+�,#��3��W�ٸ����Ok˭�g/�H��>Q�!�N�v�Ə�w��ψ��2��A�N�㻩���h�~�2��k����O� �2�xϙQ�Ƕ����Ca� $�� �B�w���X1�O�O�$�!�����6��<���<o�Ҭt���6��
��g�ފʡq�j���74�93��x����~g3t���Q�&��Z_WW�Ͻ��浶J�"Q\j?M��� w��/|X�Ŷ����7Ր�����48��[�U��!�S�r;\�yJ���:����v����4)������!��A)ISM{�����h3�� 8�!I��R�7�S���h��!0���Fl�W�������h��3��Hr����ɰ��i�o%ك�Χ���'��������V͒�+?Fy�S�{�qo��3@t�X�7�H�����s���A���t�����hCj%/un����oRщ���mF~�U���Gl-W����&����jJ���-��.�z "��v�vuή����Og�ܑV|�4��W6 zɱ$�|������YeE�����o���Վ^�t:۴�M`\����B��C*}q�6fq45/R|QM����#Նxh�P_q���U�&��,;EaE���+~�ҳo��8�PmC��*��H�֬���\$lA{d�MP7X�5�Үх�K5\�'c��������2;<��@4�~ȆA<�m�їb@�K�IWf��bpH.b~bb��s��D��#@�I��p5#{_ȃ
�Fk@������ú�����K�&�:F���U��Y������h(/���S���	!5��֩��Qޫ1�������4QGl%p~d�^]���_s��GʂIF�G�B�d�������x�P�7g�����/2g�E1p��:>%nVV''@��U���F�֬dv�|��*Q�?��&?g%HS
l0	Y�q<�۹�4��q�x|�k��T>�ݕQ{�į�1�<����8"^�o��f>N���	���!8����4�@���!L<D:Soё���'r,R�;�X��{�����4��"���[����8 ��:��^����қ��~����`J�h�"ꍳ��(�,iZ���f�k��u���0���!Bp���[�Ȫƥ�d�u�Lp�@���mu���7x�@��R��]�cC�4���%��μ�A�}�&�K�7bꅦ!����*������ =$���/�]�ϞV5�C�lKQ�{|������mK4b
�ːݿ�(��-@2�˚�\/���j�[�X���0��F��P���k@�'�o��	�j��� ��Y�J��/���.����"k� �?��Ӣ�V���%�\[d1��Am��o��yJRu˸�V�KT��S����oW�V�#����??"֒��g+|ЪG�Jj܏3�~����]nB>d�U��S��Z,j�=ɲ���>���*Ҟ�x��)�U`������2:��"�쟗T.�^&^8��i�=q��: �
����c�! �Q�3dt,m#2��v�l�"&�N��PP��C� ��=4���cev�CX�+n�W�5�Qr#4\�.2��M��l�r,�����=�.��s���6��E��C5������p��z���W%*���)�ǥ��C�\�"{�$a��'j��M^T޶���\��O�Jي��#�gM��f�!�p,/J��T��9��x�pؓ
�>���U�wP!d�D,�X��KE,Z�߫h��9.O � g��i���Q��麻g��t��Hg�rУ6{�N0�-���wwQڊS��_t��M0���7��&ٱ�LȪ�TgH��=&�3���;&��ŵ�z@���=A���2�B�앖�ͷX�4}i��>Q�y((�<I�g�t���`����Is�\���l1[f�#W93�I;ZD.3~�;�����G��P�����
XȀ�o��9ф�P�󚼼�8@6w����m�����!Ebݰn���hQ�{&��&*�)�/rdy�1����]gr]ɨ	9a]>������"��S��aL��}.��!�'VQPͣ�"�T`ޗ��C�V�e#���;M!k�;�$dq�l�;e{a��/���17 �5�P���_2ͧC�?��>Z�-ݩ�JEͶ������{kxEoB��?��\ � �����8�~�v�bIz5*�Ѻ"�x��=!�Ju����f�cw���Z
��� �ۗ�7Ɔ�:�WFN�ҡ��n`��zA�	Y��nz��=��h�\�${bˁ`@��ܱ��Y˱#�4�l�(��,�m4g��C�+�e?u�U ޫH��I�l-�Z+L]n�m�q]�V+�{�$�鎀ni
/�r(����������zf��h��״�1P&�t]���?��fDBC�>�thؙ6=��Jb�S�%�����nxD	�-�H�@}���5��%����G��/��!1�/�J��G9���)؎��_D+ե|0��՚���z�)!Q�]A���7��%�`�e��xex<�鹫�� �=��aAB&��ƥyL��:5���*�==׭�d��]%�iq�42&��q�]��E���W��"a�2'��5���żJ5S����}��S׮g��y����g\��O�a~�է�L�C��|��JE�&�L�J
��R��������y�`��*'ʜ��5I:tI^��6SB�o"z�a��=�"�+���F�F%d0�����gb$�˶�~k4M�%�A�T�/��,_%BC� �������w��<Ǉ\<�t?dw�O4��|i��*���`y2\!�f�zS�0B0��L]_p�}�;�����XI*�'��X�[i_,�$w��d������1x�"�$=)f�h����}mgW,�;��A_k����1!�E�N�贾K
�3w|�5v�\���[ڐ�v� C���iR�Y��~�Jl)���ыߊq��=�g�x��Ƣ�*����s�f�&s�ݕ_��rȠ� ׾����Bk$=���l/�N�1�^z��cD!�>0�@��*��0Z��W����3=�	ƍ���·p������=�������.�3�����N�Dk�%
�|��E�b���g��Lu��6�H�7��вA(=�4!i�"���4]�������A>�[ms*p�c}=���75�|�̇^N	�U�����q6����z���k��vˬ�H��^+�ဆ���+�57�?�=֖4bj�۟sey��|w�=��e� Z"t�%`�-s��WO����+��Z�@a��O�U#�d7���vt���em��z�r����!Aք
�ѭ��Z�qw�"�J��Y�t��	���`i{D3���W�̺f����!�߻SL��i�$o%1Yr����=���7r�$�I��\�k3�J���PGP#F\j!�O��e�


�Zk�V��B���|2������1}�:ۺ��k�������HW$���~��OUnf��.���I̮�]SL���(��� T��[Ӆt��U^�1sf��u|4����n�h
\����ٔM�����*`!Hە��=HT�	��`��'��~#�uHnh�%\Zb�:�]�fDw��hn%˲�����z�)�̑O�������'�Ǉ��s�K��kj���x�2�z¾�	Z�VufX}pqE'H�e3����\Wh\�ı�:�O~�7Y�7CH�r�O`:���*��6�_o6�l�y �p�F� mD�w�u��g�WC+:�	򣍓�
�*�'�q�cwW���ׯb!5�XR��7�7T�p������3��	�)��w4x\;�#�����C"�����()3�зj��H^�$��l�v�ʨ�ގ
����	<�����n3�貵Tǥ:
�g�͑�G��Sb�^�F?f�?Z}7�V���	p�c&eE���8&��I�������*[i-�fwܾ�:Ȑ8j��9~G:�)��mpK�;�x>�d�g�3�2N��o��gR��҂#-G߲�d��d��}\�ňH��JKL�qX~Z�jEJ��9������7��3��7q�<�u���4os�<_�!J���jqΝSF�)/�.�Sb)`2į~R��VP�'�c�8Q�I�iwh>��� �ܕ�=Wx8�����$�F���y�t5x�������3EW��rz��2G\�71mr���Ɇ��jЖ1�΢�Y�g���w6v�v�*o�;]�� �b� �/�k�7!����%bQBy%�L�e��aU?i�G<�i�Z�#i�uAD[Q�(��ϋ�4���Q`�?��_�����ys_T����Ѹ������#�]�/`��s��=.�(���q?#H�Q>�S�/F(�N�heVW�ۦl�)~yX���\�҈�lC����ۈ�ˊ_��'��fIMӾ2�I����Y<��:/k�h$��ڍ��ӔC�z?;o���<k�_OE�6jaVQL�Ά�͡�J^���ߓ�ѹD�=��,�Ɩ�M�?WE�r��}��)��y9��I��H���Y� �ߡ��p��`�H�����5��30�x%�F^$X���^+�L��4� �4�Y<`�87'��)/y]�xG�������~K�"�����)��in���=z�u�	e����X䳧�CӾ��L���ᎂ�[lΥ� �U��2���Y�3`����EV�g'���h�y�e#RB�d!td<��mYb�{��Vú�G��Ur��U�ID^JvU�B�{�є��lV{ENbAAC��e�X��TS=FG�,�q���Ӄ���=Z^�IUi�(T��W��zG�o�$�	�cL�fN�o���3�W���dl?-,���BƲ�	�H ۩,~9���90���OH���H��CiM_m�gz�ĺjL�).������f��o�G(�BOJ[RU���|�ɑ�p�
G�{=���xmq��C�����f>i'Q���8�{�����\,�uQ�b}�ɻ�f.�$�-�B�DUi8�;�K$8ię��w��/<̗;a{��/O��9&OM��S��"oz�8D����!����E9w�I"X�T���W��!:�eL�R��Dq���jg�~T�1���7#/�w��
�F���OP���&i`�43�*��B|�V,��|*���SO"�T�6i�eB����A��2�e�`� ��
B�Ȏx��M���Y����|�/��:� ��ӕ���$/�wK��)-�۔�����LƄ�:�s�F\A8��ł0��=Z�m����_�MC �i�E�:Ť��$j��ɰ~C(5��W�
F��q*E��9�O
�{a<��s�_ᄼ_�A���C��)�ߎ��y��������K���?�3.�Զ�e�OBy�w������\�fU<�Z�=e�j/�k0�Is�F���'+��&@>�&}����?��Ē)���H֜��f{/&p��L�*��R�n�[]95�C�C�օT���_�*����(aҬK��2��c����*�|���q_��|$�.KĒ�yY�i���Y���MW<>i��A8�HJ�[$ lL�k�sѭF���21��N���Z�~�YwW�J�|V�×�P64 � A}���Fw�����	mnNtX'���|��^!���`����NԸ�h&�i<����bC�mJ�@ئ�� $O���s�$������''��I0���JX%c����~S�j�B0ۿ�GO���c�U.��*a���E����(h߫F�"�F��������u��l"uz��ұ�83�h�
��{t����kh��N�ݧ�s���s��d��/�`R�7��\k�\�<�c^up_��9�]��=�O��fq���ݴ�:�ں�٘��#�>\�B�@a�Xk��u5f��~{�sY<hv�⊌���nT�q{�z�иZ&Y�|�g˕��f�%�*�g�l�LX�.��@R��_G��m=h�?FV�ʸ6���ՐT@!^| v��t^���T�v���+V��FH��L�[�K�����:*Q6���G2�N.�uG"���c@Es�7y��M�
j��،�)d?�S3(��pe����sk�N^IpY��8��پ����n����N�m���G
���͆
�������-H~?�h�=�7sj˵(32#v@tϳn�����JL25։V�����y� �l��2Q�Vp3��+�K��q�;�x���x׍��������h�v��n��H/�����;��:rq��t�``�,���Ũ^.C=r��_o%�����x�67i��>��ۅ~��\^�)=/�q�`�HÚۈ�5����.���p�l*s��EF�m7�O��v���.'�~���+�����{����ɢ��&HO>��[�5��T��F���V�z)(�m��!�hLY�ؒ�j����Y�s)��������Տ$����d��Ť�
��̋3�_r&c4�\�-�����G756� ڄ��&�������b��4c;j6�<,Hl��c��B�$�7��-ZE�i�w4�e�&ץ�e����T��h����	�R��>�7�����z'�֣��no�t����W����y��}G���'�X�{��&�������* ׼~j<��gE��a���Au��V�?��`��1��w~���[,B�=��7r&���F���F������Z��U&��/CC���~�u@	����_/�N�������J�AJ���.ZX����Q�^��j�ܖ7nv���
M>��7	���q�K��K��B�:�W,U~��=S��33<����yi��{{T����a?��6�qcKd'��ezf7jqkwt�e:x$�-�R7 �؍����Yz��{i8 -���u%^�;�@���O�迀��icQ+���ɯ�����$���V"în��y��v��\�}�8�ړ�<����9��AQ��>%���g�X֝�	��XS�}��>�7��G�]�^	@-��8�:'(��d��@�T�x�D�h���XpC�`��l�%jQ�=�V��%���f�E��)RXu	z%���,�]%�v#��Z�un�Ks�eZH�����Ņa2����9��D��� �1��5�_�h�b(�߾�A����1"�3f��	`�(�g�S[����#�������fY�AH
5Lg�"+��B� ���Y٢\�X6�M��ɾ^�������B�<)C}E8A��O@Qt�S'�6�U��e���zV)te4]nxu,ʗ�j��bꂡ��7�{[�H��^Y*w/��Au�<��=�J�`�8��i����͝+!��Mю��
|Q:��MT>�T܄!��"'ض�?�Dvd�{�n7\i���Z^8�2��۩�����Ǫ�Uqy�'Z'^�w7�4��V5h�d\��4q�D�,���i@t2W��,
�2�Z��w�@���+��M�帷����ta�>�O�
� �]f��:g1�v��ҁ�K ,[%E����Ƀ���6�c7"��@���M6�����/���vK�4�geT�� l�����П�T���׼���ɋ2Z���˚����������4\��
+���2S��4F<�[�>�6B:��E� ���1��&)�(t�,����G췳t�"�Z�bV�RRt�,����N�������r��t
'}�^�f��v� �ZN�ȑ���I\���~b�<�YO{��@E]g��l������ ���ƫ�;#��@�ذR0#nl����#+b!�j�I�A�=	u�GY��=�+|�g��u����=瑛xk.�B\�d��V���x��	����Âّ���eG�Z�ރ[��/a�W!���ɞ#�,u&	��A�.��1�|y��v�Ԃ-�)�"xt��t�.4��i_�s�ҫiy:���!.��\c���h#��wG>K�p�'m"yn9h�/SO<���ڌ70�͝hic.A� NNШBo�
�f+B�4�M�y&���J�5���,Sg��Sb[�[���}H�i��3V��#855�
B��3�g�"��u��&��`x���r�Q��:�w�ĳ�_�=��u���7�X��-�Ȟ�XN�0�"pw�ur��?G�ƫ��r� ���y�t�?����@_�w��B�M�Z!d��X�pP�BS���[����e��y0�1��� ��n�% �e�*�ܨq��� �%@>��P&��why�9�r3Z�����U��&��K��ƣʬ�'W#0���;kL��V��!����v�&�q8[%_���Ӹ�> ���կ?����.�R��{%)X��>&s C��������u"�p��ذ���U��p�܅�(mcJaN�+(�68W�J��h���~Ehy����t�Y�\��Z�2JGIu�@�R�-Њ�8�0q9�OXOѵP���Z�b��rՎ�,9�*�. �Tq'��Of�h��	~�����,rT���w�+&8���R������h�����_��#�F�?��Ɯ�^*��m	�����@�Jǹ���l���f$j[o`nI3���k2vu_z��,ܱ�[��/�(��Wt��&)��R�����l_��"|Q��C�2�C~�~'�R����W��/|7�q2�2�筝�Ɨ'�F�}})�sn��n6lޗ�u��ni��(>��_��{~	_�}�/=�{hx�	fT� qav�%n0Z���|:�@~Mv_oE�4���C�,��I�bt	|'?�6��@�BH���C��E�¶�|Y��N>�8%_%�G�Q$�ztu4d�e���H��dvZ���䍫�ЏZ��Oy��������_c��za2i��'��մ����y�s�H��>�!��Y&TTˊ�2n���|̗e�"[r(�pn
���d>l1Um�]5~��'W��(�LQA*��^SU�4xD���ѝֹu։�)Qϝ�S+���k�x�����x�W63	p����t���/d�o+�pH�0��Wx����?�a&c$[46:�Vj��+�׭�Q��_	�b���ϓ+�kP���t�XGWY�.lq���澖w<�;���Y��uL
r����w(�K��}�j6���>�\���B$��&"���ס3��5�a��ή)ߙ��K(Jj*�@���&No�l~�H�/�陹(�5��Q�#)sF���K��X7���w��?ؼ#�ڢ�יՅ�{u�ht�R����x��0�w�7����s6LЫ������Q& (�kJ'����C����z�.Z$^�[>Yp[��DN �؊:�5Y#��ʓ9E��q4I�R���� ]�F��Zz�3�d��%+h���t��ړ̷l)��K8��������ڮ��.ZY�0��$���~���St�V9+Қ��|�%��x�O�Q��s��,L[1�k���m���%��%s�-�`�@z"퀜�AkF�H1�A��-�C�cP�.�a�a��n�b�31�hA�,��>�t��1pB�
@�gҘ��40�}��<)�(R��=�X0��V���cE� t&��Er�t��q�Z��8J��g�2�iq��8�d(�Xj{�t'$�9�+[j�:<3țwq�$��6v��"��F~��w*�=�4�0`��z���7��:��n�!?[�'G'rhZ��?��T�5@�dފ
^�:��g-��_�gNE^2/��'�7WCl�0u5��xQ�<�-�� ��M�à�9��m�p�uaq�NEku�B'a�iuL��v\��iϛ�A�w�T��xen��#��I�	�4J����eϡ���עQv�ł�Ã'�+��@{�;�q�|�NrH)[��'��=Qƭ��q�2l��[l��
��;m��z@��� �7��>��C�	t<� bB��$��2���N����55P�d9�����9[fb'!M�-���A�)�㰲ͦ4R6I��ἡ�[A��xy��I��|ȥ�D�Б�Y���Cas�r��oL�Ђ�bt'	Mp����h�'�2RR��t{�L�h!`���`�/��y��5u@�p��y�ZX@Wo7z�4K`]��]����$�e���$ᬲP4k�&��H�^�!(WA�J
�Ru�P ���7k����R*�~
��/��4M�b�(c�t�ͳ��<�u�򐌲�<=��ؐ_Ei=r#�.�єO$L�.c�ÐU]��̿��͓�T��X��vo:H7�}��"!.����K�-�.��"<6']���ŉ��et����OK2Z�[����̵�;R ��
Cy��g��m�E��'��?�k8�j żwgzF�p;`E�k6�!�:cl��DC�PЖ��ڼ	�P��au�����.�٩#Y#���;��4�M�,�m0K����ߕ2�G|}��$�Mbr��;�{�Ǖ��y"�����ڡ1܈qr��4*\ߎ2���Ĉ銳W� �?�=KR�ɛ|�^n�g�W(Щǀ�����P�ϧ	�\XCj�>ë*FRx��~�ʞ�7Xd��FE�D@�B%�]hpkN�5S~]��`��u l��{�X����p^�\�%{��f�ȅ�����=��lO|z�:��i_G/&����ѕn^s@�UU ����nOcF������1��ӳN�	�^z�SuY��g�Q�������͙���^��,���K�g;���(��c�_���RsjE�;I��#��'���6�t���<�������]�=D��m�U��H���p$m������i���<_��B
�K��܌���XG!���������as�*���"�Z*��\�V� .˶|��!�w\e/�zK�N���> FU5���$�^�Vπn~����~gUtB�8^SMM���y	�6�L�1Z�F��nd�a<��ݙ]���Yщe:�|S:��%�s�{�λD�:[�N���~^�C�-t�u��dk�U.����W� t�v����XJ�H(M�\c^�3L滭�@PiË��`�jq�[3<��ϛ�*W�����_��k�@X�&�?��3��£�mC~2L��N��ذI죰�=�$$-�����p_+����7�	,�ӽ�a	R����G�y�waT4���<)0	�g5Fm��x��2�Y+9\�]/��J��Ω�h)%�Vѧ�K,jx��o^��k(�A�BQ�D��lB�y@��*	3�U���Y}��?YU�����.6U�G�:1<����m$�=��`�*]Q���+P���V��O�)HW�:�ا������r��7eʠ���:Pr%�@��|$�pV٘��C��ݼ3(!{�l��	N�u���sS�W�=�q5F��d�(�_KJ}��Q���UF�D�UNS��}۞�)�f�_/HP y+�\����"��@:\4\���H�T#UJ-
:h���dr7yg���H��*��R����??�Ɍ0e#p�%�0����sq�� ��1rw�!�`���4�Hڶj�E Mi�s�Xl�S��ݡ�F���Eܞ�ז������ik�@B赗A�X�|;�Y㠜xEH "4�,��l��b	/�;���8���ش��V�H}}~�(J(����s�(f5����]�¹#��Ű�'ڹCx8R�5'Z�+i�7q�gY~n���sϿ(�kZBMa�;ą�gԶ3�J�2�5��Oz��Q0���\ �	5(���q]M�
#����V���R=���NI2��@�^�;IH��8˱�����t�`��D�F�]�Q>�!+�xL���wE04�7P���'{"���R�'���KQWc#�6L��P~�:(�q��`X#�"�$}��R�����*N���W�ڃ�x2hH�d��GMxQ}���oǼ�8�ތ.����-�O�Ho��W�bee�'��~�M2��4�UT@�Ӊ�<y�̱��o�BVT�
�؉)z@ǟ52�,i�D��$�82�iُ�}.��m�� W"��C�{S�!b�Ğ�� cx�4�����g4�/_��/�ڼYDM���\��M:��D7O�f������aU5�s��[�Qw�_��t՘�J�m��de�CҴ@�*h(��쌌�q��_A��c��B�J���h�C���|��H���$������{�^?�
��#lu��l�Ì�5V�g��FR��&>yrT-��p�{{�47�c���_i����Ny��mڹ��t����Ѩ�pP�'vefd��4�P<q&�L]2�n�Ew���G��;n�4�ˍZ,_R��D���t�-Kϲ�@YN3�軺:��Ƙ��:j�q�%�9wV�Oe� k��מo��Q���]D:E�����1 !�H
E�+�(��/ �������%��7�L�l��)�m�w^ܣ��\�-%O��#�Bbi��4p��w�xB�&�4-�x�Kۉ��0z�����-�D$�{���g� ���ߨ��:Y�7Ai��4�B�,ˆ?��v�Ӆ���/p5�֒���גcx�2�ӦgD%N�p��ȥS\�3w7	����~����s��wVM����q����皤D��6����.8�����k�����X�-E5p)��_�,���5� �D��)&-݁���֒�f�_�l<��u��H�	0L�~�(k#6��ܶ�pdq�l�h_v	��Q����!<߷q,� E?5b�z���{�Z�ɩn��̤,�(�yz4��iF�F�.����sm�3�[�SA�ۤ� 6��p��֎*4)l�<��^3�i��Q8(�b�P/-�z�t~�CnN�}��W���xJ��FT֡ 
e���H�قA�E���t��0��=5(¬e�ᅷЍr�Sr�9v�\#2��+�7,�U�I�@��?�����F�y�oĘ�5���X�u߬n�5�Uq/W�����Q׺�G�����+h�!&*`�A�+hN���,6eU�޻ށl����%��*xo$�Z�Г�*k��!g�����me?xv�Pϕ��UĔ ��=k6/������/BR�s��ɄC7h�������z�r�URW����"lU�WJ���� Hq)i���r�>��N���`*�>J���m�e�(�4~Z\��W)$���@��Z����`t�=q�����؟�q���(s΃�r)����:Ƥ�kE7�(M�L�����)n�L0�&-+��t�O�GZ!h��Թ���5�=^�8�n�+��r�#'�	1m�x.e�����H6	בX�z=*�e��N<�a�Xa�H���&fA]!��a���x��7�W^ 2�$ �L4TO���lOo~����k5wۦ��m�uTԋ��~Tт�؄(5��{���?��A���oĝ�b��A��o�w0r^��!�|#{�����;���F�� �XVY��Հ<SwC��a�>7����������,G6i�K��$:��"V���,����(~��b�l@g�C)��ҶA�þ.�U�ZQ�K�~�M��+ZO	+?�k"�&8�������n!߽g�0��ͅ�}'��'Qa&a�Rw��?(���%ݟ�X�ֳ��>�}�

����v�i0ȑ�t�.j]~wTu���Y�����E�l`%L��+������3��T��X�<��=�A���2�l⠧�V	=�C<*���QK�N)�%b�-\C÷��V�H�S����iUq�`7��ס��L0M7dB��U��Y�7{</R����Da�����(�l�������d
p�RK��u/�|� ���>���g�w+m7Z�l�Dѿ!І�+؄�����/xp�l=
��vU�A�g��:C��~����3uS���H]����=��t~_�/�G~��~-���,D�P�k��R"���@X�SD��J��AP2��}�3�ʂ�i��6��hu`�ܽ�>�q`��:/*��%"dw��΀�q�5�����@��"�	`w��=���b��1�=R^C��QJ[��U�qaYjK�KR��Uv3���A�Bi����/��#�On����ȱs|D����h���B|��Rpߏ8����p.���|�]�T�q�gr�czM��]���"qP����tg�0�w��gg�6Fn>8��sl�F�{C#i��{�#���|��L�i�_�C(�|���\��RFT�X��y1�~_Q1�)*������ސ��m�� ��_�U�����1Rš�Z7�k-��Q9��I-�OSEFl�qa+��tXo�1�"v�Q6��ZX-k��=����/ғ��Y#�-��'YK����h�Qz�n��i�-����|��������O�5$x2���d�};>g3뱛��9\+m_�"���x�a���Y�<� T���بS �쫇��:f���}�7�_oQ���&mvk��W2�ag�|�곙��|.�F+ؖ,
~Ҫ*�٤�:�'�E��y� �h�l�ρ� Q��jZ�;x����h������9��^3ZQ��7E�[~����>Pn��o!��֡�/2�1`�v����!��ϙO��j��[,���4C���rP����77[�O�L��%ۿ�I�oi�u<�9Ǣn��6�Nf��mm(���P���ڱ�Vm��eq��f�R�-��t� ��������O��"&U�0.��P�\G(����&9ӷa�N=�
��2��� b�}�m;��r����PC�1_��؜ظ[���v��AB@��^n��ɲ�/�Z����̖&���v{#ɾ}�ws����/t�A'�{�q�����v�~��ܕ�x�
F�旺A�k$���Y�J�\��@*��o�A�k����w�����U�����:d�(O�G����#�OD��Z�����"j������j�\��;q��]����N}��y`;�3�`f��9�����(u����2p��{ ��<�I�z���Чv�E�7���_��#.j�H�x@e�v�G��R�s�pZA�`b1솋N�ê0=0�7<YR���>Eո�?7J%z�X8+%�P�AЄ��@�J�����sO7vLc��<�*��j��.���=�P��P"�Ӊq�o���E/�mN�>bc����JSG�B�������fi��$'��m�>�I�SQrqkuH���.��UA���ۍ3��ל̼�9����mFL#��M��@+[��D���LF��=���$퇑��@��IB������ FW$;*��Ǖ��I._/io��r��+|	 ɞ���PG3�wVtS�UAcu�pF]Sv��6o�������JAX���>����1118���_mDP�ۄ��O����w@	2W�r�5�7�5�0j �����W#31�6�i�Pl���$mw,��S&�Ӏ��Y�������gh�j<�6s?���rF ��qi�A�}8����k����?kp�B��ay���K�k�N!	�F:S�2�}<�M��.��E9؊�4�rF��u!t�ك�u�F+o���)%��6�+�G�������n�Yr�v}�ߗ��;F�swRr���dT�LVm�Е�����c+�C�����㼓�#��G ��+��3̈́��Y�A����	���h[:XSpX%[���&>�������q'���y�l��x^h]��)|����VKǨK��L�՗F�r���w��Y*(��:?k�=�#��6���v�{���.L���f��l��� �$��i�~V\쯨������j��*�Q�Z�TX]��4��p7��p���oM�L�c�
DG�)��ٳDӤʠRg�o�@���Ǒ�:)�m�Fi���\�O��1p�6LV�U�����ꎱM���4b����f���3���u���l���3l$x��V�'rU���4�=MKJ��8��"22���h�p�F��S�۽
��z���.��σ���sgX��������@�{F>�`0�:��<�CYȿRH����V��=�T���r��[��_�d|mMR�3�m�c��-�.Mw���t�!X����,�{u���fs�i�6�.�GD�R���<1�k�ur��J�{�@Wf�d-bi蘲�n;z���]����[M��DE��V�o/��bث���ՒM��e�O2�߱�t�#�����=����>`�[b��
üm���t�'(��b�\k,�Q�K�=��� ���.���w�@5��{�C���. Ӂ(A�� ��^���Z��>q��,JH�?P��弜���x�s��~�y���6�{"��ӈ�� ��+e?��Xr�ӄj]��nJ��!�9Ɨ��f"�����R����W��g�Oө=�V�ȦK���O$�e����B���^W�z����y��\�O���� ��g ���G!� s���{�&����.
!���q��K(^.�����+�ފ+�[䗝��s z�(Q���\���j��GE�}n�!p����V��QR���k�h�Ղ�f��Q3�O�'�߻.�m�
Jt��9�-��z�u�n@�(k�U�rI��E��}�=�]><U�����H�N;ʭ�Pʰ�7��Uj>~��r#K��ޞ��Gr�"M֜�G��^�7Bهl�;���i��[�!��̓C�c�f�h�{#/��"V�.J���y ��$7��U��?�J� �3ɅDr)���C�.������j~��H}'� '����S"��n��6g�q�}�ʐ"�~�V(Щ�rdщ�����y�����U�W18~5����{�OӗR
��Y�e�N��ɹBߛl��X`j���_�1�(5ML�>%��f�3��DM��2�;8t<�,�Q���]�
�f�����z�S�Y�F��z�s$��H���z�K'!3A��E���B�	���ﰤ�X7g����\��]���O�"��蹯�k�Y o�ŧXQ�E%>K��JP�9�Gq�+��Z�����P�b���9��]y����#�p�}������Mu���&%O��e�7�@��~��Q�P��v8)�U��8e��VNi!�����4�ͬ��Z ��t��2o{|P����ѳ@%^1��4ʊ��l�NK!��=NR�^�C,oٿ~�*��	���2�ݕ����C`3gq��kTt7����z��E`c�T	��Ֆu�]��1!K`i�%�OgJ�ծ�?��.?������S�����@�~�V_|���t���;s�X�cl�l�^_�s&�,^�h�+��[��O��!1����	�%��:d*�R���������N���k�@ڿ�ͧFc������J7�D���^I>#���5R�G�q�'����ض�uq�U-�L�P���>H�/���#�u�ο���2�؝�d�&�A�[W:c��n��Q�>2�����a�v/](%H��a#�_(xk�~�8�?`a�ϑ��T�6�7�;��)��5�4�s��=_�-!\�vF�o{Yp�O��	@���x}`k�.d]���B��1��?���~��s���9BY�ݵ��������@;��Xo
�I�-]ӊ�����S4�Ld�f�̐�6w��p��u걟�N/H\�U7�3�s�lˎa��y��3 6�9o����R��8�MY��=����� �=U�t�Y�Ґd8�ЛFT��y8�Uy����ۭ{j�	�n�P'y�K&J�[�jQ��z�%F�*�a�&��Us��L�%�5�B�o���XA���M�b�F�q��j��*�@.�q~�}CzI0
5I"�٩r�s��8���G����H˵|2�[��"2���S���٫�F�ԄS��d}���ڋR��m���Ќ��MDM|�)�6TN.��� ,�W�# �O��|���*�uБ����fPd"�( ���1{ut�� `�������J���V� $�ka�����k%��O0b&TT�G �������GG@ n���C�XV�S�� X*x���ZKQ�]W�4e�IU0N�{�E��p*���z.�h�!�-��^[�`�sT^¸�M^�	�u�K�}b�H�9F��x��G,����*Z�R1�g�M���%�c����]��C�DG�gЗP��3ůǤDØg:��R�X���@�K�i�0gSvD^�U�p���]�'�-���q�V��z+�v�\��3<��1�-����V\ʱ}*��Az�A�; �b�� ߅�,�Q)V��sD�au����Mh��ɗ_}�d�h�Nk�D�R�z����Y�ą�3_�/�a�U��{��δ��|+�X�SE�D�
�M~�]���ХIը�	]�����>��It�[]Nr2��9�R�)(Ý�c�#< ^�P���K���cw��j�� 	U9�H�4��K��\S�.&�q�Ŵ0���m�J=�V3��@7=�D���l����.�sw�Fz��;x���z�I��5�C��PL\��ټ[�7����s�W���XH�ݗ W�{�P�3ϋ�gS��>#��I��E���ڌF�m�L�~U����Zj%}�c�*�в��b�� ����������u-��ϕ��π�Q#1hs�kL"m�poA���M���Zĥ!�U�[�v<է�;� �t�����n�f����@:�!������	ڋ��Mw��������DiAk��q�k<��Y�`����&ff4�F�[�&�9뤏$B"�6!�����㍵�og�3����h'�*@Ɲ�(&%��8�Ȕ��(��~@o3��`�Q��گ��g��I	 '���0��T/ʥ]����x�
`	���5���/�'p�8�ғ�DrýI9�݄�7�uo���X�)K��ڽ8��u;}�Ml8x�Rm��B����$%xj5�c�!#	�$�#�GY�L^�)���:�_���&'�f��U�?�	~�b �