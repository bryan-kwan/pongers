// top_level.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module top_level (
		output wire        audio_out_writeresponsevalid_n, //              audio_out.writeresponsevalid_n
		input  wire        clk_clk,                        //                    clk.clk
		input  wire [3:0]  gpio_export,                    //                   gpio.export
		output wire [12:0] memory_addr,                    //                 memory.addr
		output wire [1:0]  memory_ba,                      //                       .ba
		output wire        memory_cas_n,                   //                       .cas_n
		output wire        memory_cke,                     //                       .cke
		output wire        memory_cs_n,                    //                       .cs_n
		inout  wire [15:0] memory_dq,                      //                       .dq
		output wire [1:0]  memory_dqm,                     //                       .dqm
		output wire        memory_ras_n,                   //                       .ras_n
		output wire        memory_we_n,                    //                       .we_n
		output wire        sdram_clk_clk,                  //              sdram_clk.clk
		input  wire        spi_master_MISO,                //             spi_master.MISO
		output wire        spi_master_MOSI,                //                       .MOSI
		output wire        spi_master_SCLK,                //                       .SCLK
		output wire        spi_master_SS_n,                //                       .SS_n
		output wire        spi_slave_MISO,                 //              spi_slave.MISO
		input  wire        spi_slave_MOSI,                 //                       .MOSI
		input  wire        spi_slave_SCLK,                 //                       .SCLK
		input  wire        spi_slave_SS_n,                 //                       .SS_n
		input  wire [7:0]  sw_external_connection_export,  // sw_external_connection.export
		output wire        vga_conduit_CLK,                //            vga_conduit.CLK
		output wire        vga_conduit_HS,                 //                       .HS
		output wire        vga_conduit_VS,                 //                       .VS
		output wire        vga_conduit_BLANK,              //                       .BLANK
		output wire        vga_conduit_SYNC,               //                       .SYNC
		output wire [3:0]  vga_conduit_R,                  //                       .R
		output wire [3:0]  vga_conduit_G,                  //                       .G
		output wire [3:0]  vga_conduit_B                   //                       .B
	);

	wire         video_alpha_blender_0_avalon_blended_source_valid;                                        // video_alpha_blender_0:output_valid -> video_dual_clock_buffer_0:stream_in_valid
	wire  [29:0] video_alpha_blender_0_avalon_blended_source_data;                                         // video_alpha_blender_0:output_data -> video_dual_clock_buffer_0:stream_in_data
	wire         video_alpha_blender_0_avalon_blended_source_ready;                                        // video_dual_clock_buffer_0:stream_in_ready -> video_alpha_blender_0:output_ready
	wire         video_alpha_blender_0_avalon_blended_source_startofpacket;                                // video_alpha_blender_0:output_startofpacket -> video_dual_clock_buffer_0:stream_in_startofpacket
	wire         video_alpha_blender_0_avalon_blended_source_endofpacket;                                  // video_alpha_blender_0:output_endofpacket -> video_dual_clock_buffer_0:stream_in_endofpacket
	wire         video_character_buffer_with_dma_0_avalon_char_source_valid;                               // video_character_buffer_with_dma_0:stream_valid -> video_alpha_blender_0:foreground_valid
	wire  [39:0] video_character_buffer_with_dma_0_avalon_char_source_data;                                // video_character_buffer_with_dma_0:stream_data -> video_alpha_blender_0:foreground_data
	wire         video_character_buffer_with_dma_0_avalon_char_source_ready;                               // video_alpha_blender_0:foreground_ready -> video_character_buffer_with_dma_0:stream_ready
	wire         video_character_buffer_with_dma_0_avalon_char_source_startofpacket;                       // video_character_buffer_with_dma_0:stream_startofpacket -> video_alpha_blender_0:foreground_startofpacket
	wire         video_character_buffer_with_dma_0_avalon_char_source_endofpacket;                         // video_character_buffer_with_dma_0:stream_endofpacket -> video_alpha_blender_0:foreground_endofpacket
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_valid;                                  // video_dual_clock_buffer_0:stream_out_valid -> video_vga_controller_0:valid
	wire  [29:0] video_dual_clock_buffer_0_avalon_dc_buffer_source_data;                                   // video_dual_clock_buffer_0:stream_out_data -> video_vga_controller_0:data
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_ready;                                  // video_vga_controller_0:ready -> video_dual_clock_buffer_0:stream_out_ready
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket;                          // video_dual_clock_buffer_0:stream_out_startofpacket -> video_vga_controller_0:startofpacket
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket;                            // video_dual_clock_buffer_0:stream_out_endofpacket -> video_vga_controller_0:endofpacket
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_valid;                                       // video_pixel_buffer_dma_0:stream_valid -> video_rgb_resampler_0:stream_in_valid
	wire  [15:0] video_pixel_buffer_dma_0_avalon_pixel_source_data;                                        // video_pixel_buffer_dma_0:stream_data -> video_rgb_resampler_0:stream_in_data
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_ready;                                       // video_rgb_resampler_0:stream_in_ready -> video_pixel_buffer_dma_0:stream_ready
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket;                               // video_pixel_buffer_dma_0:stream_startofpacket -> video_rgb_resampler_0:stream_in_startofpacket
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket;                                 // video_pixel_buffer_dma_0:stream_endofpacket -> video_rgb_resampler_0:stream_in_endofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_valid;                                            // video_rgb_resampler_0:stream_out_valid -> video_scaler_0:stream_in_valid
	wire  [29:0] video_rgb_resampler_0_avalon_rgb_source_data;                                             // video_rgb_resampler_0:stream_out_data -> video_scaler_0:stream_in_data
	wire         video_rgb_resampler_0_avalon_rgb_source_ready;                                            // video_scaler_0:stream_in_ready -> video_rgb_resampler_0:stream_out_ready
	wire         video_rgb_resampler_0_avalon_rgb_source_startofpacket;                                    // video_rgb_resampler_0:stream_out_startofpacket -> video_scaler_0:stream_in_startofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_endofpacket;                                      // video_rgb_resampler_0:stream_out_endofpacket -> video_scaler_0:stream_in_endofpacket
	wire         altpll_0_c0_clk;                                                                          // altpll_0:c0 -> [audio_module_0:clock25, rst_controller_002:clk, video_dual_clock_buffer_0:clk_stream_out, video_vga_controller_0:clk]
	wire         top_level_debug_reset_request_reset;                                                      // top_level:debug_reset_request -> [mm_interconnect_0:spi_0_reset_reset_bridge_in_reset_reset, rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_001:reset_in1, rst_controller_002:reset_in0, spi_0:reset_n, spi_1:reset_n]
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest;                             // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest -> video_pixel_buffer_dma_0:master_waitrequest
	wire  [15:0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata;                                // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata -> video_pixel_buffer_dma_0:master_readdata
	wire  [31:0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_address;                                 // video_pixel_buffer_dma_0:master_address -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_address
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_read;                                    // video_pixel_buffer_dma_0:master_read -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_read
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid;                           // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid -> video_pixel_buffer_dma_0:master_readdatavalid
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock;                                    // video_pixel_buffer_dma_0:master_arbiterlock -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock
	wire  [31:0] top_level_data_master_readdata;                                                           // mm_interconnect_0:top_level_data_master_readdata -> top_level:d_readdata
	wire         top_level_data_master_waitrequest;                                                        // mm_interconnect_0:top_level_data_master_waitrequest -> top_level:d_waitrequest
	wire         top_level_data_master_debugaccess;                                                        // top_level:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:top_level_data_master_debugaccess
	wire  [27:0] top_level_data_master_address;                                                            // top_level:d_address -> mm_interconnect_0:top_level_data_master_address
	wire   [3:0] top_level_data_master_byteenable;                                                         // top_level:d_byteenable -> mm_interconnect_0:top_level_data_master_byteenable
	wire         top_level_data_master_read;                                                               // top_level:d_read -> mm_interconnect_0:top_level_data_master_read
	wire         top_level_data_master_write;                                                              // top_level:d_write -> mm_interconnect_0:top_level_data_master_write
	wire  [31:0] top_level_data_master_writedata;                                                          // top_level:d_writedata -> mm_interconnect_0:top_level_data_master_writedata
	wire  [31:0] top_level_instruction_master_readdata;                                                    // mm_interconnect_0:top_level_instruction_master_readdata -> top_level:i_readdata
	wire         top_level_instruction_master_waitrequest;                                                 // mm_interconnect_0:top_level_instruction_master_waitrequest -> top_level:i_waitrequest
	wire  [27:0] top_level_instruction_master_address;                                                     // top_level:i_address -> mm_interconnect_0:top_level_instruction_master_address
	wire         top_level_instruction_master_read;                                                        // top_level:i_read -> mm_interconnect_0:top_level_instruction_master_read
	wire         mm_interconnect_0_new_sdram_controller_0_s1_chipselect;                                   // mm_interconnect_0:new_sdram_controller_0_s1_chipselect -> new_sdram_controller_0:az_cs
	wire  [15:0] mm_interconnect_0_new_sdram_controller_0_s1_readdata;                                     // new_sdram_controller_0:za_data -> mm_interconnect_0:new_sdram_controller_0_s1_readdata
	wire         mm_interconnect_0_new_sdram_controller_0_s1_waitrequest;                                  // new_sdram_controller_0:za_waitrequest -> mm_interconnect_0:new_sdram_controller_0_s1_waitrequest
	wire  [24:0] mm_interconnect_0_new_sdram_controller_0_s1_address;                                      // mm_interconnect_0:new_sdram_controller_0_s1_address -> new_sdram_controller_0:az_addr
	wire         mm_interconnect_0_new_sdram_controller_0_s1_read;                                         // mm_interconnect_0:new_sdram_controller_0_s1_read -> new_sdram_controller_0:az_rd_n
	wire   [1:0] mm_interconnect_0_new_sdram_controller_0_s1_byteenable;                                   // mm_interconnect_0:new_sdram_controller_0_s1_byteenable -> new_sdram_controller_0:az_be_n
	wire         mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid;                                // new_sdram_controller_0:za_valid -> mm_interconnect_0:new_sdram_controller_0_s1_readdatavalid
	wire         mm_interconnect_0_new_sdram_controller_0_s1_write;                                        // mm_interconnect_0:new_sdram_controller_0_s1_write -> new_sdram_controller_0:az_wr_n
	wire  [15:0] mm_interconnect_0_new_sdram_controller_0_s1_writedata;                                    // mm_interconnect_0:new_sdram_controller_0_s1_writedata -> new_sdram_controller_0:az_data
	wire  [31:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata;                 // video_pixel_buffer_dma_0:slave_readdata -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_readdata
	wire   [1:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address;                  // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_address -> video_pixel_buffer_dma_0:slave_address
	wire         mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read;                     // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_read -> video_pixel_buffer_dma_0:slave_read
	wire   [3:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable;               // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_byteenable -> video_pixel_buffer_dma_0:slave_byteenable
	wire         mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write;                    // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_write -> video_pixel_buffer_dma_0:slave_write
	wire  [31:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata;                // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_writedata -> video_pixel_buffer_dma_0:slave_writedata
	wire  [31:0] mm_interconnect_0_top_level_debug_mem_slave_readdata;                                     // top_level:debug_mem_slave_readdata -> mm_interconnect_0:top_level_debug_mem_slave_readdata
	wire         mm_interconnect_0_top_level_debug_mem_slave_waitrequest;                                  // top_level:debug_mem_slave_waitrequest -> mm_interconnect_0:top_level_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_top_level_debug_mem_slave_debugaccess;                                  // mm_interconnect_0:top_level_debug_mem_slave_debugaccess -> top_level:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_top_level_debug_mem_slave_address;                                      // mm_interconnect_0:top_level_debug_mem_slave_address -> top_level:debug_mem_slave_address
	wire         mm_interconnect_0_top_level_debug_mem_slave_read;                                         // mm_interconnect_0:top_level_debug_mem_slave_read -> top_level:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_top_level_debug_mem_slave_byteenable;                                   // mm_interconnect_0:top_level_debug_mem_slave_byteenable -> top_level:debug_mem_slave_byteenable
	wire         mm_interconnect_0_top_level_debug_mem_slave_write;                                        // mm_interconnect_0:top_level_debug_mem_slave_write -> top_level:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_top_level_debug_mem_slave_writedata;                                    // mm_interconnect_0:top_level_debug_mem_slave_writedata -> top_level:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                                         // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                                           // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory2_0_s1_address;                                            // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                                         // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                                              // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                                          // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                                              // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_timer_0_s1_chipselect;                                                  // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                                                    // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                                                     // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                                                       // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                                                   // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect;  // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect -> video_character_buffer_with_dma_0:buf_chipselect
	wire   [7:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata;    // video_character_buffer_with_dma_0:buf_readdata -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest; // video_character_buffer_with_dma_0:buf_waitrequest -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest
	wire  [12:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address;     // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_address -> video_character_buffer_with_dma_0:buf_address
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read;        // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_read -> video_character_buffer_with_dma_0:buf_read
	wire   [0:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable;  // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable -> video_character_buffer_with_dma_0:buf_byteenable
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write;       // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_write -> video_character_buffer_with_dma_0:buf_write
	wire   [7:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata;   // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata -> video_character_buffer_with_dma_0:buf_writedata
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect; // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect -> video_character_buffer_with_dma_0:ctrl_chipselect
	wire  [31:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata;   // video_character_buffer_with_dma_0:ctrl_readdata -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_readdata
	wire   [0:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address;    // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_address -> video_character_buffer_with_dma_0:ctrl_address
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read;       // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_read -> video_character_buffer_with_dma_0:ctrl_read
	wire   [3:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable; // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable -> video_character_buffer_with_dma_0:ctrl_byteenable
	wire         mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write;      // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_write -> video_character_buffer_with_dma_0:ctrl_write
	wire  [31:0] mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata;  // mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_writedata -> video_character_buffer_with_dma_0:ctrl_writedata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;                               // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;                                 // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;                              // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;                                  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;                                     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;                                    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;                                // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_audio_module_0_avalon_slave_0_1_readdata;                               // audio_module_0:readdata -> mm_interconnect_0:audio_module_0_avalon_slave_0_1_readdata
	wire         mm_interconnect_0_audio_module_0_avalon_slave_0_1_read;                                   // mm_interconnect_0:audio_module_0_avalon_slave_0_1_read -> audio_module_0:read
	wire         mm_interconnect_0_audio_module_0_avalon_slave_0_1_write;                                  // mm_interconnect_0:audio_module_0_avalon_slave_0_1_write -> audio_module_0:write
	wire  [31:0] mm_interconnect_0_audio_module_0_avalon_slave_0_1_writedata;                              // mm_interconnect_0:audio_module_0_avalon_slave_0_1_writedata -> audio_module_0:writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;                                    // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;                                     // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;                                            // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;                                             // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                                                // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                                               // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;                                           // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire         mm_interconnect_0_sw_s1_chipselect;                                                       // mm_interconnect_0:sw_s1_chipselect -> sw:chipselect
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                                                         // sw:readdata -> mm_interconnect_0:sw_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                                                          // mm_interconnect_0:sw_s1_address -> sw:address
	wire         mm_interconnect_0_sw_s1_write;                                                            // mm_interconnect_0:sw_s1_write -> sw:write_n
	wire  [31:0] mm_interconnect_0_sw_s1_writedata;                                                        // mm_interconnect_0:sw_s1_writedata -> sw:writedata
	wire         mm_interconnect_0_gpio_s1_chipselect;                                                     // mm_interconnect_0:GPIO_s1_chipselect -> GPIO:chipselect
	wire  [31:0] mm_interconnect_0_gpio_s1_readdata;                                                       // GPIO:readdata -> mm_interconnect_0:GPIO_s1_readdata
	wire   [1:0] mm_interconnect_0_gpio_s1_address;                                                        // mm_interconnect_0:GPIO_s1_address -> GPIO:address
	wire         mm_interconnect_0_gpio_s1_write;                                                          // mm_interconnect_0:GPIO_s1_write -> GPIO:write_n
	wire  [31:0] mm_interconnect_0_gpio_s1_writedata;                                                      // mm_interconnect_0:GPIO_s1_writedata -> GPIO:writedata
	wire         mm_interconnect_0_spi_0_spi_control_port_chipselect;                                      // mm_interconnect_0:spi_0_spi_control_port_chipselect -> spi_0:spi_select
	wire  [15:0] mm_interconnect_0_spi_0_spi_control_port_readdata;                                        // spi_0:data_to_cpu -> mm_interconnect_0:spi_0_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_0_spi_control_port_address;                                         // mm_interconnect_0:spi_0_spi_control_port_address -> spi_0:mem_addr
	wire         mm_interconnect_0_spi_0_spi_control_port_read;                                            // mm_interconnect_0:spi_0_spi_control_port_read -> spi_0:read_n
	wire         mm_interconnect_0_spi_0_spi_control_port_write;                                           // mm_interconnect_0:spi_0_spi_control_port_write -> spi_0:write_n
	wire  [15:0] mm_interconnect_0_spi_0_spi_control_port_writedata;                                       // mm_interconnect_0:spi_0_spi_control_port_writedata -> spi_0:data_from_cpu
	wire         mm_interconnect_0_spi_1_spi_control_port_chipselect;                                      // mm_interconnect_0:spi_1_spi_control_port_chipselect -> spi_1:spi_select
	wire  [15:0] mm_interconnect_0_spi_1_spi_control_port_readdata;                                        // spi_1:data_to_cpu -> mm_interconnect_0:spi_1_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_1_spi_control_port_address;                                         // mm_interconnect_0:spi_1_spi_control_port_address -> spi_1:mem_addr
	wire         mm_interconnect_0_spi_1_spi_control_port_read;                                            // mm_interconnect_0:spi_1_spi_control_port_read -> spi_1:read_n
	wire         mm_interconnect_0_spi_1_spi_control_port_write;                                           // mm_interconnect_0:spi_1_spi_control_port_write -> spi_1:write_n
	wire  [15:0] mm_interconnect_0_spi_1_spi_control_port_writedata;                                       // mm_interconnect_0:spi_1_spi_control_port_writedata -> spi_1:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                                                 // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                 // timer_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                                 // sw:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                                 // GPIO:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                                 // spi_0:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                                                 // spi_1:irq -> irq_mapper:receiver5_irq
	wire  [31:0] top_level_irq_irq;                                                                        // irq_mapper:sender_irq -> top_level:irq
	wire         video_scaler_0_avalon_scaler_source_valid;                                                // video_scaler_0:stream_out_valid -> avalon_st_adapter:in_0_valid
	wire  [29:0] video_scaler_0_avalon_scaler_source_data;                                                 // video_scaler_0:stream_out_data -> avalon_st_adapter:in_0_data
	wire         video_scaler_0_avalon_scaler_source_ready;                                                // avalon_st_adapter:in_0_ready -> video_scaler_0:stream_out_ready
	wire   [1:0] video_scaler_0_avalon_scaler_source_channel;                                              // video_scaler_0:stream_out_channel -> avalon_st_adapter:in_0_channel
	wire         video_scaler_0_avalon_scaler_source_startofpacket;                                        // video_scaler_0:stream_out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         video_scaler_0_avalon_scaler_source_endofpacket;                                          // video_scaler_0:stream_out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire         avalon_st_adapter_out_0_valid;                                                            // avalon_st_adapter:out_0_valid -> video_alpha_blender_0:background_valid
	wire  [29:0] avalon_st_adapter_out_0_data;                                                             // avalon_st_adapter:out_0_data -> video_alpha_blender_0:background_data
	wire         avalon_st_adapter_out_0_ready;                                                            // video_alpha_blender_0:background_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                                                    // avalon_st_adapter:out_0_startofpacket -> video_alpha_blender_0:background_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                                                      // avalon_st_adapter:out_0_endofpacket -> video_alpha_blender_0:background_endofpacket
	wire         rst_controller_reset_out_reset;                                                           // rst_controller:reset_out -> [GPIO:reset_n, altpll_0:reset, audio_module_0:reset_n, avalon_st_adapter:in_rst_0_reset, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:video_pixel_buffer_dma_0_reset_reset_bridge_in_reset_reset, new_sdram_controller_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, sw:reset_n, sysid_qsys_0:reset_n, timer_0:reset_n, top_level:reset_n, video_dual_clock_buffer_0:reset_stream_in, video_pixel_buffer_dma_0:reset, video_rgb_resampler_0:reset, video_scaler_0:reset]
	wire         rst_controller_reset_out_reset_req;                                                       // rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in, top_level:reset_req]
	wire         rst_controller_001_reset_out_reset;                                                       // rst_controller_001:reset_out -> [mm_interconnect_0:video_character_buffer_with_dma_0_reset_reset_bridge_in_reset_reset, video_alpha_blender_0:reset, video_character_buffer_with_dma_0:reset]
	wire         rst_controller_002_reset_out_reset;                                                       // rst_controller_002:reset_out -> [video_dual_clock_buffer_0:reset_stream_out, video_vga_controller_0:reset]

	top_level_GPIO gpio (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_gpio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpio_s1_readdata),   //                    .readdata
		.in_port    (gpio_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)              //                 irq.irq
	);

	top_level_altpll_0 altpll_0 (
		.clk                (clk_clk),                                        //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset),                 // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_0_c0_clk),                                //                    c0.clk
		.c1                 (),                                               //                    c1.clk
		.locked             (),                                               //        locked_conduit.export
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.c2                 (),                                               //           (terminated)
		.c3                 (),                                               //           (terminated)
		.c4                 (),                                               //           (terminated)
		.areset             (1'b0),                                           //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (3'b000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	audio_avalon_interface audio_module_0 (
		.reset_n   (~rst_controller_reset_out_reset),                             //      clock_reset.reset_n
		.speaker   (audio_out_writeresponsevalid_n),                              //      conduit_end.writeresponsevalid_n
		.clock25   (altpll_0_c0_clk),                                             //    clock_sink_25.clk
		.clock50   (clk_clk),                                                     //    clock_sink_50.clk
		.writedata (mm_interconnect_0_audio_module_0_avalon_slave_0_1_writedata), // avalon_slave_0_1.writedata
		.write     (mm_interconnect_0_audio_module_0_avalon_slave_0_1_write),     //                 .write
		.read      (mm_interconnect_0_audio_module_0_avalon_slave_0_1_read),      //                 .read
		.readdata  (mm_interconnect_0_audio_module_0_avalon_slave_0_1_readdata)   //                 .readdata
	);

	top_level_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	top_level_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (clk_clk),                                                   //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                           // reset.reset_n
		.az_addr        (mm_interconnect_0_new_sdram_controller_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_new_sdram_controller_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_new_sdram_controller_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_new_sdram_controller_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_new_sdram_controller_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_new_sdram_controller_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (memory_addr),                                               //  wire.export
		.zs_ba          (memory_ba),                                                 //      .export
		.zs_cas_n       (memory_cas_n),                                              //      .export
		.zs_cke         (memory_cke),                                                //      .export
		.zs_cs_n        (memory_cs_n),                                               //      .export
		.zs_dq          (memory_dq),                                                 //      .export
		.zs_dqm         (memory_dqm),                                                //      .export
		.zs_ras_n       (memory_ras_n),                                              //      .export
		.zs_we_n        (memory_we_n)                                                //      .export
	);

	top_level_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	top_level_spi_0 spi_0 (
		.clk           (clk_clk),                                             //              clk.clk
		.reset_n       (~top_level_debug_reset_request_reset),                //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_0_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_0_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_0_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_0_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_0_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_0_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver4_irq),                            //              irq.irq
		.MISO          (spi_slave_MISO),                                      //         external.export
		.MOSI          (spi_slave_MOSI),                                      //                 .export
		.SCLK          (spi_slave_SCLK),                                      //                 .export
		.SS_n          (spi_slave_SS_n)                                       //                 .export
	);

	top_level_spi_1 spi_1 (
		.clk           (clk_clk),                                             //              clk.clk
		.reset_n       (~top_level_debug_reset_request_reset),                //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_1_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_1_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_1_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_1_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_1_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_1_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver5_irq),                            //              irq.irq
		.MISO          (spi_master_MISO),                                     //         external.export
		.MOSI          (spi_master_MOSI),                                     //                 .export
		.SCLK          (spi_master_SCLK),                                     //                 .export
		.SS_n          (spi_master_SS_n)                                      //                 .export
	);

	top_level_sw sw (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_sw_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sw_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sw_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sw_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sw_s1_readdata),   //                    .readdata
		.in_port    (sw_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver2_irq)            //                 irq.irq
	);

	top_level_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	top_level_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	top_level_top_level top_level (
		.clk                                 (clk_clk),                                                 //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                         //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                      //                          .reset_req
		.d_address                           (top_level_data_master_address),                           //               data_master.address
		.d_byteenable                        (top_level_data_master_byteenable),                        //                          .byteenable
		.d_read                              (top_level_data_master_read),                              //                          .read
		.d_readdata                          (top_level_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (top_level_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (top_level_data_master_write),                             //                          .write
		.d_writedata                         (top_level_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (top_level_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (top_level_instruction_master_address),                    //        instruction_master.address
		.i_read                              (top_level_instruction_master_read),                       //                          .read
		.i_readdata                          (top_level_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (top_level_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (top_level_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (top_level_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_top_level_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_top_level_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_top_level_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_top_level_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_top_level_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_top_level_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_top_level_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_top_level_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                         // custom_instruction_master.readra
	);

	top_level_video_alpha_blender_0 video_alpha_blender_0 (
		.clk                      (clk_clk),                                                            //                    clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                 //                  reset.reset
		.foreground_data          (video_character_buffer_with_dma_0_avalon_char_source_data),          // avalon_foreground_sink.data
		.foreground_startofpacket (video_character_buffer_with_dma_0_avalon_char_source_startofpacket), //                       .startofpacket
		.foreground_endofpacket   (video_character_buffer_with_dma_0_avalon_char_source_endofpacket),   //                       .endofpacket
		.foreground_valid         (video_character_buffer_with_dma_0_avalon_char_source_valid),         //                       .valid
		.foreground_ready         (video_character_buffer_with_dma_0_avalon_char_source_ready),         //                       .ready
		.background_data          (avalon_st_adapter_out_0_data),                                       // avalon_background_sink.data
		.background_startofpacket (avalon_st_adapter_out_0_startofpacket),                              //                       .startofpacket
		.background_endofpacket   (avalon_st_adapter_out_0_endofpacket),                                //                       .endofpacket
		.background_valid         (avalon_st_adapter_out_0_valid),                                      //                       .valid
		.background_ready         (avalon_st_adapter_out_0_ready),                                      //                       .ready
		.output_ready             (video_alpha_blender_0_avalon_blended_source_ready),                  //  avalon_blended_source.ready
		.output_data              (video_alpha_blender_0_avalon_blended_source_data),                   //                       .data
		.output_startofpacket     (video_alpha_blender_0_avalon_blended_source_startofpacket),          //                       .startofpacket
		.output_endofpacket       (video_alpha_blender_0_avalon_blended_source_endofpacket),            //                       .endofpacket
		.output_valid             (video_alpha_blender_0_avalon_blended_source_valid)                   //                       .valid
	);

	top_level_video_character_buffer_with_dma_0 video_character_buffer_with_dma_0 (
		.clk                  (clk_clk),                                                                                  //                       clk.clk
		.reset                (rst_controller_001_reset_out_reset),                                                       //                     reset.reset
		.ctrl_address         (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable), //                          .byteenable
		.ctrl_chipselect      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect), //                          .chipselect
		.ctrl_read            (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read),       //                          .read
		.ctrl_write           (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write),      //                          .write
		.ctrl_writedata       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata),  //                          .writedata
		.ctrl_readdata        (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata),   //                          .readdata
		.buf_byteenable       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect),  //                          .chipselect
		.buf_read             (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read),        //                          .read
		.buf_write            (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write),       //                          .write
		.buf_writedata        (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata),   //                          .writedata
		.buf_readdata         (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata),    //                          .readdata
		.buf_waitrequest      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest), //                          .waitrequest
		.buf_address          (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address),     //                          .address
		.stream_ready         (video_character_buffer_with_dma_0_avalon_char_source_ready),                               //        avalon_char_source.ready
		.stream_startofpacket (video_character_buffer_with_dma_0_avalon_char_source_startofpacket),                       //                          .startofpacket
		.stream_endofpacket   (video_character_buffer_with_dma_0_avalon_char_source_endofpacket),                         //                          .endofpacket
		.stream_valid         (video_character_buffer_with_dma_0_avalon_char_source_valid),                               //                          .valid
		.stream_data          (video_character_buffer_with_dma_0_avalon_char_source_data)                                 //                          .data
	);

	top_level_video_dual_clock_buffer_0 video_dual_clock_buffer_0 (
		.clk_stream_in            (clk_clk),                                                         //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                                  //         reset_stream_in.reset
		.clk_stream_out           (altpll_0_c0_clk),                                                 //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_002_reset_out_reset),                              //        reset_stream_out.reset
		.stream_in_ready          (video_alpha_blender_0_avalon_blended_source_ready),               //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (video_alpha_blender_0_avalon_blended_source_startofpacket),       //                        .startofpacket
		.stream_in_endofpacket    (video_alpha_blender_0_avalon_blended_source_endofpacket),         //                        .endofpacket
		.stream_in_valid          (video_alpha_blender_0_avalon_blended_source_valid),               //                        .valid
		.stream_in_data           (video_alpha_blender_0_avalon_blended_source_data),                //                        .data
		.stream_out_ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data)           //                        .data
	);

	top_level_video_pixel_buffer_dma_0 video_pixel_buffer_dma_0 (
		.clk                  (clk_clk),                                                                    //                     clk.clk
		.reset                (rst_controller_reset_out_reset),                                             //                   reset.reset
		.master_readdatavalid (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid),             // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest),               //                        .waitrequest
		.master_address       (video_pixel_buffer_dma_0_avalon_pixel_dma_master_address),                   //                        .address
		.master_arbiterlock   (video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock),                      //                        .lock
		.master_read          (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read),                      //                        .read
		.master_readdata      (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata),                  //                        .readdata
		.slave_address        (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address),    //    avalon_control_slave.address
		.slave_byteenable     (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable), //                        .byteenable
		.slave_read           (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read),       //                        .read
		.slave_write          (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write),      //                        .write
		.slave_writedata      (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata),  //                        .writedata
		.slave_readdata       (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata),   //                        .readdata
		.stream_ready         (video_pixel_buffer_dma_0_avalon_pixel_source_ready),                         //     avalon_pixel_source.ready
		.stream_startofpacket (video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket),                 //                        .startofpacket
		.stream_endofpacket   (video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket),                   //                        .endofpacket
		.stream_valid         (video_pixel_buffer_dma_0_avalon_pixel_source_valid),                         //                        .valid
		.stream_data          (video_pixel_buffer_dma_0_avalon_pixel_source_data)                           //                        .data
	);

	top_level_video_rgb_resampler_0 video_rgb_resampler_0 (
		.clk                      (clk_clk),                                                    //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                             //             reset.reset
		.stream_in_startofpacket  (video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (video_pixel_buffer_dma_0_avalon_pixel_source_valid),         //                  .valid
		.stream_in_ready          (video_pixel_buffer_dma_0_avalon_pixel_source_ready),         //                  .ready
		.stream_in_data           (video_pixel_buffer_dma_0_avalon_pixel_source_data),          //                  .data
		.stream_out_ready         (video_rgb_resampler_0_avalon_rgb_source_ready),              // avalon_rgb_source.ready
		.stream_out_startofpacket (video_rgb_resampler_0_avalon_rgb_source_startofpacket),      //                  .startofpacket
		.stream_out_endofpacket   (video_rgb_resampler_0_avalon_rgb_source_endofpacket),        //                  .endofpacket
		.stream_out_valid         (video_rgb_resampler_0_avalon_rgb_source_valid),              //                  .valid
		.stream_out_data          (video_rgb_resampler_0_avalon_rgb_source_data)                //                  .data
	);

	top_level_video_scaler_0 video_scaler_0 (
		.clk                      (clk_clk),                                               //                  clk.clk
		.reset                    (rst_controller_reset_out_reset),                        //                reset.reset
		.stream_in_startofpacket  (video_rgb_resampler_0_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (video_rgb_resampler_0_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (video_rgb_resampler_0_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (video_rgb_resampler_0_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (video_rgb_resampler_0_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (video_scaler_0_avalon_scaler_source_ready),             // avalon_scaler_source.ready
		.stream_out_startofpacket (video_scaler_0_avalon_scaler_source_startofpacket),     //                     .startofpacket
		.stream_out_endofpacket   (video_scaler_0_avalon_scaler_source_endofpacket),       //                     .endofpacket
		.stream_out_valid         (video_scaler_0_avalon_scaler_source_valid),             //                     .valid
		.stream_out_data          (video_scaler_0_avalon_scaler_source_data),              //                     .data
		.stream_out_channel       (video_scaler_0_avalon_scaler_source_channel)            //                     .channel
	);

	top_level_video_vga_controller_0 video_vga_controller_0 (
		.clk           (altpll_0_c0_clk),                                                 //                clk.clk
		.reset         (rst_controller_002_reset_out_reset),                              //              reset.reset
		.data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_conduit_CLK),                                                 // external_interface.export
		.VGA_HS        (vga_conduit_HS),                                                  //                   .export
		.VGA_VS        (vga_conduit_VS),                                                  //                   .export
		.VGA_BLANK     (vga_conduit_BLANK),                                               //                   .export
		.VGA_SYNC      (vga_conduit_SYNC),                                                //                   .export
		.VGA_R         (vga_conduit_R),                                                   //                   .export
		.VGA_G         (vga_conduit_G),                                                   //                   .export
		.VGA_B         (vga_conduit_B)                                                    //                   .export
	);

	top_level_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                                          (clk_clk),                                                                                  //                                                     clk_0_clk.clk
		.spi_0_reset_reset_bridge_in_reset_reset                                (top_level_debug_reset_request_reset),                                                      //                             spi_0_reset_reset_bridge_in_reset.reset
		.video_character_buffer_with_dma_0_reset_reset_bridge_in_reset_reset    (rst_controller_001_reset_out_reset),                                                       // video_character_buffer_with_dma_0_reset_reset_bridge_in_reset.reset
		.video_pixel_buffer_dma_0_reset_reset_bridge_in_reset_reset             (rst_controller_reset_out_reset),                                                           //          video_pixel_buffer_dma_0_reset_reset_bridge_in_reset.reset
		.top_level_data_master_address                                          (top_level_data_master_address),                                                            //                                         top_level_data_master.address
		.top_level_data_master_waitrequest                                      (top_level_data_master_waitrequest),                                                        //                                                              .waitrequest
		.top_level_data_master_byteenable                                       (top_level_data_master_byteenable),                                                         //                                                              .byteenable
		.top_level_data_master_read                                             (top_level_data_master_read),                                                               //                                                              .read
		.top_level_data_master_readdata                                         (top_level_data_master_readdata),                                                           //                                                              .readdata
		.top_level_data_master_write                                            (top_level_data_master_write),                                                              //                                                              .write
		.top_level_data_master_writedata                                        (top_level_data_master_writedata),                                                          //                                                              .writedata
		.top_level_data_master_debugaccess                                      (top_level_data_master_debugaccess),                                                        //                                                              .debugaccess
		.top_level_instruction_master_address                                   (top_level_instruction_master_address),                                                     //                                  top_level_instruction_master.address
		.top_level_instruction_master_waitrequest                               (top_level_instruction_master_waitrequest),                                                 //                                                              .waitrequest
		.top_level_instruction_master_read                                      (top_level_instruction_master_read),                                                        //                                                              .read
		.top_level_instruction_master_readdata                                  (top_level_instruction_master_readdata),                                                    //                                                              .readdata
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_address               (video_pixel_buffer_dma_0_avalon_pixel_dma_master_address),                                 //              video_pixel_buffer_dma_0_avalon_pixel_dma_master.address
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest           (video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest),                             //                                                              .waitrequest
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_read                  (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read),                                    //                                                              .read
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata              (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata),                                //                                                              .readdata
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid         (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid),                           //                                                              .readdatavalid
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock                  (video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock),                                    //                                                              .lock
		.altpll_0_pll_slave_address                                             (mm_interconnect_0_altpll_0_pll_slave_address),                                             //                                            altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                               (mm_interconnect_0_altpll_0_pll_slave_write),                                               //                                                              .write
		.altpll_0_pll_slave_read                                                (mm_interconnect_0_altpll_0_pll_slave_read),                                                //                                                              .read
		.altpll_0_pll_slave_readdata                                            (mm_interconnect_0_altpll_0_pll_slave_readdata),                                            //                                                              .readdata
		.altpll_0_pll_slave_writedata                                           (mm_interconnect_0_altpll_0_pll_slave_writedata),                                           //                                                              .writedata
		.audio_module_0_avalon_slave_0_1_write                                  (mm_interconnect_0_audio_module_0_avalon_slave_0_1_write),                                  //                               audio_module_0_avalon_slave_0_1.write
		.audio_module_0_avalon_slave_0_1_read                                   (mm_interconnect_0_audio_module_0_avalon_slave_0_1_read),                                   //                                                              .read
		.audio_module_0_avalon_slave_0_1_readdata                               (mm_interconnect_0_audio_module_0_avalon_slave_0_1_readdata),                               //                                                              .readdata
		.audio_module_0_avalon_slave_0_1_writedata                              (mm_interconnect_0_audio_module_0_avalon_slave_0_1_writedata),                              //                                                              .writedata
		.GPIO_s1_address                                                        (mm_interconnect_0_gpio_s1_address),                                                        //                                                       GPIO_s1.address
		.GPIO_s1_write                                                          (mm_interconnect_0_gpio_s1_write),                                                          //                                                              .write
		.GPIO_s1_readdata                                                       (mm_interconnect_0_gpio_s1_readdata),                                                       //                                                              .readdata
		.GPIO_s1_writedata                                                      (mm_interconnect_0_gpio_s1_writedata),                                                      //                                                              .writedata
		.GPIO_s1_chipselect                                                     (mm_interconnect_0_gpio_s1_chipselect),                                                     //                                                              .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),                                  //                                 jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),                                    //                                                              .write
		.jtag_uart_0_avalon_jtag_slave_read                                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),                                     //                                                              .read
		.jtag_uart_0_avalon_jtag_slave_readdata                                 (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),                                 //                                                              .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),                                //                                                              .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),                              //                                                              .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),                               //                                                              .chipselect
		.new_sdram_controller_0_s1_address                                      (mm_interconnect_0_new_sdram_controller_0_s1_address),                                      //                                     new_sdram_controller_0_s1.address
		.new_sdram_controller_0_s1_write                                        (mm_interconnect_0_new_sdram_controller_0_s1_write),                                        //                                                              .write
		.new_sdram_controller_0_s1_read                                         (mm_interconnect_0_new_sdram_controller_0_s1_read),                                         //                                                              .read
		.new_sdram_controller_0_s1_readdata                                     (mm_interconnect_0_new_sdram_controller_0_s1_readdata),                                     //                                                              .readdata
		.new_sdram_controller_0_s1_writedata                                    (mm_interconnect_0_new_sdram_controller_0_s1_writedata),                                    //                                                              .writedata
		.new_sdram_controller_0_s1_byteenable                                   (mm_interconnect_0_new_sdram_controller_0_s1_byteenable),                                   //                                                              .byteenable
		.new_sdram_controller_0_s1_readdatavalid                                (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid),                                //                                                              .readdatavalid
		.new_sdram_controller_0_s1_waitrequest                                  (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),                                  //                                                              .waitrequest
		.new_sdram_controller_0_s1_chipselect                                   (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),                                   //                                                              .chipselect
		.onchip_memory2_0_s1_address                                            (mm_interconnect_0_onchip_memory2_0_s1_address),                                            //                                           onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                              (mm_interconnect_0_onchip_memory2_0_s1_write),                                              //                                                              .write
		.onchip_memory2_0_s1_readdata                                           (mm_interconnect_0_onchip_memory2_0_s1_readdata),                                           //                                                              .readdata
		.onchip_memory2_0_s1_writedata                                          (mm_interconnect_0_onchip_memory2_0_s1_writedata),                                          //                                                              .writedata
		.onchip_memory2_0_s1_byteenable                                         (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                                         //                                                              .byteenable
		.onchip_memory2_0_s1_chipselect                                         (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                                         //                                                              .chipselect
		.onchip_memory2_0_s1_clken                                              (mm_interconnect_0_onchip_memory2_0_s1_clken),                                              //                                                              .clken
		.spi_0_spi_control_port_address                                         (mm_interconnect_0_spi_0_spi_control_port_address),                                         //                                        spi_0_spi_control_port.address
		.spi_0_spi_control_port_write                                           (mm_interconnect_0_spi_0_spi_control_port_write),                                           //                                                              .write
		.spi_0_spi_control_port_read                                            (mm_interconnect_0_spi_0_spi_control_port_read),                                            //                                                              .read
		.spi_0_spi_control_port_readdata                                        (mm_interconnect_0_spi_0_spi_control_port_readdata),                                        //                                                              .readdata
		.spi_0_spi_control_port_writedata                                       (mm_interconnect_0_spi_0_spi_control_port_writedata),                                       //                                                              .writedata
		.spi_0_spi_control_port_chipselect                                      (mm_interconnect_0_spi_0_spi_control_port_chipselect),                                      //                                                              .chipselect
		.spi_1_spi_control_port_address                                         (mm_interconnect_0_spi_1_spi_control_port_address),                                         //                                        spi_1_spi_control_port.address
		.spi_1_spi_control_port_write                                           (mm_interconnect_0_spi_1_spi_control_port_write),                                           //                                                              .write
		.spi_1_spi_control_port_read                                            (mm_interconnect_0_spi_1_spi_control_port_read),                                            //                                                              .read
		.spi_1_spi_control_port_readdata                                        (mm_interconnect_0_spi_1_spi_control_port_readdata),                                        //                                                              .readdata
		.spi_1_spi_control_port_writedata                                       (mm_interconnect_0_spi_1_spi_control_port_writedata),                                       //                                                              .writedata
		.spi_1_spi_control_port_chipselect                                      (mm_interconnect_0_spi_1_spi_control_port_chipselect),                                      //                                                              .chipselect
		.sw_s1_address                                                          (mm_interconnect_0_sw_s1_address),                                                          //                                                         sw_s1.address
		.sw_s1_write                                                            (mm_interconnect_0_sw_s1_write),                                                            //                                                              .write
		.sw_s1_readdata                                                         (mm_interconnect_0_sw_s1_readdata),                                                         //                                                              .readdata
		.sw_s1_writedata                                                        (mm_interconnect_0_sw_s1_writedata),                                                        //                                                              .writedata
		.sw_s1_chipselect                                                       (mm_interconnect_0_sw_s1_chipselect),                                                       //                                                              .chipselect
		.sysid_qsys_0_control_slave_address                                     (mm_interconnect_0_sysid_qsys_0_control_slave_address),                                     //                                    sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                                    (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),                                    //                                                              .readdata
		.timer_0_s1_address                                                     (mm_interconnect_0_timer_0_s1_address),                                                     //                                                    timer_0_s1.address
		.timer_0_s1_write                                                       (mm_interconnect_0_timer_0_s1_write),                                                       //                                                              .write
		.timer_0_s1_readdata                                                    (mm_interconnect_0_timer_0_s1_readdata),                                                    //                                                              .readdata
		.timer_0_s1_writedata                                                   (mm_interconnect_0_timer_0_s1_writedata),                                                   //                                                              .writedata
		.timer_0_s1_chipselect                                                  (mm_interconnect_0_timer_0_s1_chipselect),                                                  //                                                              .chipselect
		.top_level_debug_mem_slave_address                                      (mm_interconnect_0_top_level_debug_mem_slave_address),                                      //                                     top_level_debug_mem_slave.address
		.top_level_debug_mem_slave_write                                        (mm_interconnect_0_top_level_debug_mem_slave_write),                                        //                                                              .write
		.top_level_debug_mem_slave_read                                         (mm_interconnect_0_top_level_debug_mem_slave_read),                                         //                                                              .read
		.top_level_debug_mem_slave_readdata                                     (mm_interconnect_0_top_level_debug_mem_slave_readdata),                                     //                                                              .readdata
		.top_level_debug_mem_slave_writedata                                    (mm_interconnect_0_top_level_debug_mem_slave_writedata),                                    //                                                              .writedata
		.top_level_debug_mem_slave_byteenable                                   (mm_interconnect_0_top_level_debug_mem_slave_byteenable),                                   //                                                              .byteenable
		.top_level_debug_mem_slave_waitrequest                                  (mm_interconnect_0_top_level_debug_mem_slave_waitrequest),                                  //                                                              .waitrequest
		.top_level_debug_mem_slave_debugaccess                                  (mm_interconnect_0_top_level_debug_mem_slave_debugaccess),                                  //                                                              .debugaccess
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_address     (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address),     //    video_character_buffer_with_dma_0_avalon_char_buffer_slave.address
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_write       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write),       //                                                              .write
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_read        (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read),        //                                                              .read
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata    (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata),    //                                                              .readdata
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata   (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata),   //                                                              .writedata
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable  (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable),  //                                                              .byteenable
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest), //                                                              .waitrequest
		.video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect  (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect),  //                                                              .chipselect
		.video_character_buffer_with_dma_0_avalon_char_control_slave_address    (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address),    //   video_character_buffer_with_dma_0_avalon_char_control_slave.address
		.video_character_buffer_with_dma_0_avalon_char_control_slave_write      (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write),      //                                                              .write
		.video_character_buffer_with_dma_0_avalon_char_control_slave_read       (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read),       //                                                              .read
		.video_character_buffer_with_dma_0_avalon_char_control_slave_readdata   (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata),   //                                                              .readdata
		.video_character_buffer_with_dma_0_avalon_char_control_slave_writedata  (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata),  //                                                              .writedata
		.video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable), //                                                              .byteenable
		.video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect (mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect), //                                                              .chipselect
		.video_pixel_buffer_dma_0_avalon_control_slave_address                  (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address),                  //                 video_pixel_buffer_dma_0_avalon_control_slave.address
		.video_pixel_buffer_dma_0_avalon_control_slave_write                    (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write),                    //                                                              .write
		.video_pixel_buffer_dma_0_avalon_control_slave_read                     (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read),                     //                                                              .read
		.video_pixel_buffer_dma_0_avalon_control_slave_readdata                 (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata),                 //                                                              .readdata
		.video_pixel_buffer_dma_0_avalon_control_slave_writedata                (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata),                //                                                              .writedata
		.video_pixel_buffer_dma_0_avalon_control_slave_byteenable               (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable)                //                                                              .byteenable
	);

	top_level_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.sender_irq    (top_level_irq_irq)               //    sender.irq
	);

	top_level_avalon_st_adapter #(
		.inBitsPerSymbol (10),
		.inUsePackets    (1),
		.inDataWidth     (30),
		.inChannelWidth  (2),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (30),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                                           // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),                    // in_rst_0.reset
		.in_0_data           (video_scaler_0_avalon_scaler_source_data),          //     in_0.data
		.in_0_valid          (video_scaler_0_avalon_scaler_source_valid),         //         .valid
		.in_0_ready          (video_scaler_0_avalon_scaler_source_ready),         //         .ready
		.in_0_startofpacket  (video_scaler_0_avalon_scaler_source_startofpacket), //         .startofpacket
		.in_0_endofpacket    (video_scaler_0_avalon_scaler_source_endofpacket),   //         .endofpacket
		.in_0_channel        (video_scaler_0_avalon_scaler_source_channel),       //         .channel
		.out_0_data          (avalon_st_adapter_out_0_data),                      //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                     //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                     //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),             //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)                //         .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (top_level_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_in1      (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (top_level_debug_reset_request_reset), // reset_in0.reset
		.reset_in1      (top_level_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (top_level_debug_reset_request_reset), // reset_in0.reset
		.clk            (altpll_0_c0_clk),                     //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_in1      (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	assign sdram_clk_clk = clk_clk;

endmodule
