��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����{hi��7	G�����|��4/���YEs��Q��H�9e���ϒ��(��t�.�?�ѩ<�Փ�<�Evj���T�����B�ݰ7� ػ�3��p�����D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�������+�%ix��;��-���y��6XM�F���
]8.�"y5��[S��I~o03�v�4�W�����x���W��>!�3�i�/�T���Q\�^u���?��bUc3�̠�"x� V�ǁ��}�0��*{7�uY�v�]�fr�$ݦ��x,q�@�?\�q*��g�����q�0��T�*��Ϭ~����pCl��>����4�s���K%�_EDi�b��}�bB���<��ٟRg���J-�7`?��x��¬�n�t��d�\�K�[[庢]߾�)ӷǏ�ӑރ�TQ���b�sq�*͘x�[O?�c ^yKH0U՝6����6�f���{D�+��n�cK��h�ߜ<l��"«e���mx��!m�~o��\$��kK���8*�M}.�>�/����������4�?�#rN�g�Gpi���v/

k����c]�]�(����&兵����GUW�*�P��5C���jcBH��D z�G��_�40�����>�^@М뀏��=eU�6���tx�m$�7���\���qI��ݫ}廈	��B���/$vTYɳ�:�T!0�D�q9Br�b�O����l�W$��c��m� _�V�qX�������z7�}�� 6�^л���	)=+6|Ng���<0�%����m��l_ah��P����% &p=r�n�%66��8�f��^���[\��1��~��7�����.Ӥ�y@�d�=V���������J�$�y�Q��:'����ɨ�8�����L-z|��z��`l���'>��pd�[jV�1ҡ.c�7xx��k�÷e�f�`�x��Q�O���;*��A���B呙/��@ҥ��;���������f �L(A�X������SU��F���T�l��S⠪y��8�Ԕ�v �#��[6�۩�ɝw��(%������t���^��k���Y&�w��ĤY�Pz���|���/+3A����\;��H��\��{�a�3Z�`�j>�E��3DY,s|� "�:��*�@��<�*��2�ywG��`x@��Rl[����@(TG��i�7㵝�p)�O��������@�xY�~��S�v�� ֚�m6�.{��)��I��	?��o��P�j��&� �ʴ�h���z���/Q)��U.ym.�լr(h���;��<ԣ��]Yt|�|V�G,���!Iq�$ަU�<0�g��U%��}#���e����64��u��}Fճ��K��1}�W��9���R68k.l[s,e�s������׹,�bal�����P��m�B���ט�{\}Wm��|h��1�-�m|��m������㯸9	�}��t�:�@9�[Zs���1�����k�2C@)�Іg�P��,���"��|(��ԑ�cY�:��Zv_YA��5���V�Xs����Hn}�q�c9���ͦ��D̑`ވ���vc+aw�)O���q�N�y>S�K�)9�2�6�-��U�n�|�b���q��|o6��;�k2fG�A�!��1�~���j
ZS���,2"��������%��,�ɊrI�~�x���~ý�c-��d1)/�oW�_P,���㝁ZV�>�6�F>UD��%���E9J�f�Qo]x=�[G�%���ï��_�)�JNl}O�^�m�v&e���zSfɒ�ڒ+V�V���EY�������q���8�"x�1K�1�������?��4KtJ��%A��������R@ɪ�������q1��$��8����ȥ��l�nP�Ġrw��+-�j��e�5�Քkze�|�'�$�
�\S�e:�C�R��7i#�-1�ac��S�4�z�F{��
2�-�1����c<���q�n+�fk�n�J�lw$|y�����ZϮ���z���-��^:B=�P.��z����<w�lφ�7Q�R����}�]bǐ�<I�2Lf'�kT��������[�|s�95
ɣ�K4։����тa�{P�&e�9/�]xT�TM�,���-�R�����!��{A��e���m�2p�~{��!=�Z��E�6J�@Q�'C��m��@%������w�qd��]�k�Ӑ>Y�2[�gtU˹�I;���g闻���֐եc��\R��ى����ɓ��ߧ)!FG�� y��F�W�+BLbob�-M�jަ�d�O�W���>;|�.��~7�j;T���4h����l�d�3:�ŉ�D>�ö��@�G�2�m��ݮQqЫk�6���b*<u���C���W�4>�lƨ��='�@��'�`*��O34�V���`�\�������Ŀ2�)z���Ƶ����
����GJt�uôk-Y����\հ�F����o<�'MVr7>Y�ջ#߶	f�f�i8��x�k�h<�!*O��ະ�X��,%�/;9_�R����䐣�8bf���]��$� �g�:<.x�5p����
����(6=W:K^���5�T��~���8����^����X��:e�YxdF��w������i';�Q��y��|+r����Ï�"N�mG�,��r��E�o��2;X�72J=��
�W�u���`�?�-]�ْ%	�.PB
ƺ`G<Y�b�xܙP8R�S��(D�9K�J%/*le�i�ȓ)�p���B7m�B;��2f���6ëZ
��`���� ���FJ���A���~��^�C��gy���/�&"�m�/omfi5�F�[��G�wb gx��s+�����ʹ8{~(B�q��)hTcݭZ��7��;����|���ӳ��;Y���~�ّ�0IF=`DGPRRp�e?��9�G_��J��%
K���4��S�h�l��I�ʋ��y�.#[�ʮ��`*A�Jw;�yZ���X,�Ir��̐I�\�a]ט��i��x�J���m|��~�og�{{
Ch�c>�����%��x�򤳘��e�5D�=�]}�������k=�w�ra�^�ª�����e�G���_n*֖!�:�N"���/p�޳��gZ�X�J��K$�U�F�ka۟��r��-XO�Ï�E���o����
q�z�M/��f�Mq9]ݷ8�.0-<)�8�4؃�ht�m��.M��ߏPqn&>�61^U�5/F��#3����f:?KP��0%nF[.���a��K�~7�fz<�/�&���
�&����kب����a7m��R�r%���?+��aKc?��^�c�����#�C�����,Vh0$������Y܃�4,���@�Ի��[/���bE_�_�fn�\Q�
�X>�+�;�lՆ�
κ��{����,�ts�$�՚3|����P�v��9����<�QF^�Da�,�7���`x�L��Bp��%��F��x�g6w�si$ݺX?D��ֵzOf�#(Q�a�	�iYN��BMZ.�23��L��¾	��62yn�i���E��=
7�I��&����${�K��I�i��O�/��<n�I�L�W�ܩ���o��?B��`��.��4�u��p����r�	 FyocV�h�t�#�"s�#���� i���̥����i���ȭ���'�h�a#qN_/k~�uק�<T�7%r�6"!	fZ�"��d�U���o����?Ȋ�M�F (,�{X�EJ?%���}��4'�S7��sQ|�I�>|ӿ�v�!|�c�����T =u�ɰlu�>ƬPͳy�|�o�±�bR5 ��Hm<6`WB<N޻�JV�F��KE�H�Vj>2gPv��0<c�MY��CA��.Y��<��h�����["�MH�c�:����&xW��9���?������|�O�lJ=����+���`��;���O�^�UHM�a�U���^�A�}$���W��|���>���-�¶'��i�Wl527��̎ŲX�a�hx6U��t'qL�s*:;��J�w��3ϥ��A���;���E�Y��ax�z��'�Ү���&�Ixl��L::�Ļ*��y�OϾ�|��%�X�cJ����V�� 6�K�*��+Pn�/c�c�ڌ��K�����Ji����� ��J�JOP]�H���S�,�����Y���S�i)NG\�N�B�&��6��l�>��+�:��� o ���¤t֖��X>\P�9�k�⅊�wuf��蠽��d��`3�^��)5!���B�+uR�Q/~�g���~��^��D�v�=��G'�}��}�%�zP�����6�ǧ�����R����,ђ_"�tA{�j�BA�_���P��&�Ո	S�sW�̓�u��$x�;��Q�ξ��Ǵ�ƹ`��%V0�}�'�SNw��:O����
/X3�I,D���wx�p�W����$P���Į�����m�Wi�n@�|�涨fg*InN���=�.�����B������9MsQ���ۥ���$u�\ �Ji����܄x������cY�~����':�BWI�����juhv7ie�M�u�n@�*�9�I!-��o�����G�L֋h{]���<���Ml�R,Y��"�sL�����p�����|kDt��ɕ%��#H�sa��|;ԇ�}5�����"�f�"����1C8���>��S(�`{�Y[��&��}ka��RԌw�:�OL��+ol3��-,@]�Q�@�:�̀m�c�D����{���d�[aܙH�_4��E���&I��$2ś�#�n��',��+���=���
�Ӕ����K#�Ģ+1��IpZ�`��v��i޾d���WU|G���^2�h�<����= ��i�R��m5��
0N��֑�|L����{��%ĽƄ�Ⴀ����/��h�nk��ǣЩ���]�KH?�h�'M�F�8PM�������O��Nb�t�[��"��c]��~�
��0������E�-���6R�.k� c���Q���3D�$K�YőWs�bH���k���ÙK��!G(`V��S�����J?j�a@�5�.+
�"Ma��[�yf%��N&"�4�U����zxC-�� �w$%��`J��q���6	T���֌�M���+��������A�5L��D������=�t*�cK�[��7H���K�v����D�YK`f��x�7�=�^��:�T�K����FQ)U8��n�(F�<4�S!;��؟�z��m[�����,���w��XsT��d��w�y��Sw���e��������y���%�/����F����o�R`_懼P��b�[g��w�I��l��v��j�����\ZS��1p���kۘ����9�eh����P����g�VPMZ���j7C9[K��uD;h�Q���D����Og���q(�/Z2���pu�_&UYr��ɢ��>ް֏<��!eDз�}����N��H�|��kN)�-_�*��R~����rΧJܨgԹШr燲�l"���!`�A܃�A �`�YN�Gn���(�֯��
�8�6b�{qً��L�Q���Lmv����5������"t�`��h�>�q���*N|�����=W�+�Ya�H�hn�V���.c������2��R?*���^+�<�*�wY���f|2�6�(�Y�:��x�2���z���δc��u�o�R��d�@�U��	8
�~�������Z�q'���2��_P�KV����S��$qܗE^�%�$��e���,j�(��v��Fx�0���1V��΁��D�j+���nĖ����,��}3��c����VO0S�zfv���B�}W[���NjwE^w
�A��0�p���-ʰ۾��@#6~�܄O��B���y�V*FSk��b�(zJ��������qM�ҡ�2�0cXY�=�n� �B)�v��E}�SUr!�X�/�]�`����R�d�pݦ2� i��15�ֺh�H̛�X%�����8�� �~�{�*���Er�����>:� ���Zl�،�\��-)���"@�(�I`�z��*�nz��`k{�(�M��O.ғ�J�L��4���kqH\�h��o"������!ERq!TI}��;����JV(?���Y,�s���5�;'&��-�&�f�)�Cy��G���xn���m`C'B-�����j�3�/�8�W�	��]�EX�t�u1Z�rj��i�ҟ�\Ŧ#�V���iӗ��Ç�BVHR[kJ|&h5qz#(.�_s���D���O����Þ��ĝ��R�FM%h��9E[	IS�J;����	��ᨓ�]ס�_+^����2�|�9O��ݔY�u�*��m��c�,�T�˖�����r7��JG�4v��ZJ��a��1�k�0� �f�O+虯;@c?������B���A�H��G1�~��q�/>��aF�B�1�X���>�4�i�w
���L S��`O0_-z�}�:A�s�{Z�O/Xn��W5s�xu�3�q�=���jɷ�ǳ��i!cF���%��HH"Q2����V�q���s�*����Lx�Ɇן��T��W�e�÷#�������+7��9�0W�%z�Y�ñ�3���IL�W�(���3�9������U�Ψ����!6l	��8-;˩&ɻ�"-,�Eý!��3��	 �W�3S������ <��귤������k����,G��1%2n5�XUXz�E�Я�qV���8�M������+rź#��~z�T�E���2(�z����z�v����T}��9��뤊@,�=�y�'U�V�c������d�[�D��Kh�՜xt����@Gx��9��w�0 ��:]�����h^�n�G�����T��$��~5���]RM�������a��2�h���'���@�h\wU`nX����{d��� B���;��:L
�(�~������^F-p�g���eM3l�+���B�i��o}v-Yo�����~Xa�9f�T�w�ZW�@đ�09�0�Y\���I��ܜ�L(� ���+L'X�ꂑ{d�ۃ�E��K�����~�:]�L?������vwz	 _�S,��,��W�+P@�8�`�Z��d}#=%I���'�k}'t�41��K]2n����&��lID0oטp0^���3�Jܭ�c(t����vk�+�~7w�ǸL*n�|���a�ˏ�Tv��� '��-GH$��v�j��[���'jd3�'V��C�w1vr�o#. ��׫���)Z�������7�Մ��0�|^:Uؗ%��ɏ�����Z�Z!���͵]��z��9*�	o���<���^��<	p�Aw����`�y�`C�3�r��~8�����C�4֔+t���dl��jn�ӯ_��I1Jө�Ս�*o�3���9I2��c��Қ�x6�X��\��A�'ʁb�x߹<�ӕ[#�b���K�O�\A�W!})}
D��\E`����3Z��;"�YX�+����-)=5��L���	h��"���zU/+��.=�1�}��qB?L�H����Ӟ͇YPf�- VR��;���u9r�+��y�Y�.��U���9±6� RH]�O��.�榇{����˞{'/���c�#Vm����|�E�փRN�I��{�~mRRIFv�HV��J�	�Y��G���NO�����ß�3�$@⩫���� �d<3�F��'9�*�T3��[�i�S3�Y����u#���9Vk���c���:+�5"���툿.����x�L[�������9����m��-c�!�n[�g����M�ݚ�4B����{g|�9�N�^~]��yp*1ʅިOZIy���b8˜�[}���&�u�L�L�4Ȯ��73��/�����N��[�0������BR\����g���x�C�&sL �jpd�@p�4�,��d�X�	���"�;E��:���cA�Î�4+�Lv�y&�V���! ��*�\s�n�V菛�ٺ*�LgŋcnEc~G�p(�0E�:t/v?�n<����ć4�`[����*��d��xZ�ղ%����2D�D8�h�%��\�ҮN��_� �D���_;P�-d�ʄ�q�;���O�}�<"<�֪Yc���d�z�F�(��>F%��X�h���6f���o��d�����݈:���鮵�G�&g��P�~j,&Z�,ހ��x �$��ȯf���x@V��s�S{�����@d#`����SYߟ�H�����i}S,��QU1@��Bj�׈���ȃ�RE���f;�����Q��4�|��m�� p"�zE�������X�Z�>迭���QN����X\��;e����8w\�6��{����t5�9oa��{�=q�,�?׊�-B�&��Z���85�o6��r�E�/�#���j�jzHW�Q��%fd�C��h�peo��Ƹ.,�LGX�������3�7/8-K��?�O@2_�ن̐#�����s�=��{���S�7��&���o��,d}liK\[�H�Y���ϤwM���+b�ͮZ�n��R��z,hPje���$=��i�N����{�- :�ɵ T�_m���YLV' �F�3��6D�����%����r�eBK�w�k[�v�)W/,6U��B	ѭ�wg��|G���9��.Q{9��yip MT懈��F%E%/߸o��E�p��jX����B��޻ws�U�mp�����H,_PVw��;{�g!���p<8��[�Jg��Vw�����(��v~*>{�
_���J<��;��.ٚ�o��sOs�r؛�h�t? I��sn�!o��*ݒ%�^!�rVm�ڎh8˅�[�A/�
 ����"���٣Ω� ΁�n�y	�y���7H��K+��/;{�ep3���^����{�f}`�d-�Q�5��%K�� �C:��~�;Nx������y�}x�6�
霆 ��3��,_[�c�	Ԁ���9Q�ȫM�}������|`΢�+|�QF�jSA蛨��^ؘa���� ��\�FI>҂"u4}��z��������8.?������C<e�����,���F�)�v�eɜvKbͳ��>k�>�[U=��?�������D�����[��7E��.I���'�<��?�������O4Vh���^A�H)Q[�b��q�X�^�%Œ[+�t�: uE���4X�g��+10���"G��5}�;�ᕽy71�ubL�I-(#�t�G"`�>Zh��ʚ>� �G���;��<�B}���\]�ԥ�6_��̯l]��?#��%���p��H�+�Z2U�΢	|Ǉ�DL�I�,�������GǶĦ�j�:=)b	��|-K�"IC����R	���I6ˎLH���L6��<�W��.���׿�bH%5�//3I��͂���>6c�a�R�7�i���h&�C床��u,@ۥ)�rw��B��F�v� �(8_�a�HC��A��i�i5��F����x^��*w���&�ɦ���.�z5��w�`%��u�n���
1�RNr���Xb��Z�y�?V�� �Pbm�������*�Mĺ�0�cgn�ws�yh�6����!�N�u:�����BGa��Y2�� �$�eD�R0���vTv�5��F(�~�]t(�c�ٴ {>Q�KV���S����b� 9��޵��S �H 5C}+x�c15T���������˶j��kڬ�C7�vESk`��b�zRVNc{�2���m�%�[Y�"���F'0���/�4�̅��Р�[. �[�;ŘK_�w��pO���[vˌ|�M�Z)�<������ŭ�A\.+� N�c
�I�����������s�*_��$��[Z/�I�${6=����E�oo$����*f5�2_u�R���m��	�S��8ӐqA��؝�wG�0�^`�*zbSL��U��W��r>G����ڂ���$\Ue,vw��\4d��&��:#o����9s�}�����$�F�JCE!\��T9=�!��:��>�#T|2���J3~��n-�8vg�(���EK�b(pTeq-�+	N�^�1��?
�����{��(/s`ς�*y�i)��Ƌ��Zpm$�ӈMg��sf�=�ƽux'��93��M���O��'T���spJ�
��t��0�7�ʎ^�l�lRL+d+��I��7���m[�ԓ�{��ȩ	�*�^��jI7f��d	�Lf��Vg�|T�>��L"�Ĩ�GHe!!
<�>��4���� /�y��\��VLc�|���` �/�D����L�)<�h�&&p5'��a��Cy�?���e�ɝ�:"��<cl�a��Gu�b�����\}0p&�na���'�K�Π�G���˧ExU� +n��R��>��x�DIn��@Y�Ӌ����ќ@�d�<��9	�GOC�����-dJ:'ۿ���:D"��6�D.�Ar*��u�����j����Xٝ��t��oJ��E����h�`y������o�����2Q-ڼ�L���84�m��d ��]Kԛ�jW@?�>�0 4�e�;^��-��������1�`�q��eO�������̋��'
g�Zao]��\b]xv�g����%rLo�X��#��֛�~?��f|�	i�n%��M4y�.���W� �����ƯF�(��Û��[��C�����M-��j�=wE��	�{���wm�:+.|�q�0j~WH�W�0<p9�L�8��F�<���	^����	W��o&��O���m��d8T�_+�.�6n�(�q1��}�<g|V��d�f=�Ά�X͂���a]R5&R��	��:h���PzzzV鸁r�����/����3�n1�S/\Є�}��'�l�HR�\�!�N\/���7M����dE*|޳
�.��U.����v�὘�1��~��/�lK��#�;����5ϾC����e��O���k�}���J;��r�qn:ZA���M/���Y8�)wg2U�%�)ǀr�5RRgc!Yۅ�l3���Y�-�w�-a�i��3��.�'s���Q��:�z~�$�a�Fʳ� FI�!a����ҠԦ��q�������3�3�DDjٴh�����G��dh�|�����tw�Q?��8��5m�ćg�`� !�2�kXJ��c�ߝZrN�uo�.m���ǿ*	�W�U��q��o�q>���
H|b��r烧X�kj!��ipj|ơ��y�b��U�翑s����ԫ�
�$�
�����u��|��Zu�mD��s�Ӝ'2�g���d�X"&x���i;5~�K�8 t�����'�dqgD�#�ɧ���2�e#nK+?�ȴ$�����.G�P'�+��/j��Y��Rm$�K�ŧ(��T^
B�*6@���/�X���mQ��g�-:��O3���bAtm�\��e�
��<��XGͫ'9�)q��n&��)�6�O��8�)'�ӧ��2�M)��$ZkdH׸�{���4�|����)�QԽ ���Ќ�ȑ���C����v�<���"w4L)NL��ͪv�#G�2�#AS��^<�ϧ�*w�� �]�<�%�Kf�b�w�-o�ЩǪ�%.�v�IO�<')TV�H��=$���Or�9�v/޳���6��ؼ�Y�|���1�����iB��C��ͫ�Ҳ��T9dB��4�Xk_��g��1 [�� ݆�<#\&����,�5z�C=eB��}�_J̥fAϦ&��I֜
��JX��?�[�ہ	�[�S���V������h4 �2�P�\\�4�s6�Z���ߦܷty�/u��	0vMY�!��$���BVeN��&
5ՂHp`,k�%�5v�4�y�o��ͩ3
tT��~U✝�;ڧ�@��d0d�E��ղ4<K7)��eJiIa_���gvʬ�6�+Ǭ5g��an���m���o�o>�p�i��sit۟׶6�YZ^�p���(KQe���R��)�Q��G�ɧJ���%��3�ㄵtM�H�Dr��F� �
F8�d�/*Xp�vZW��q�8gf%��%��>{�cUU��B�Ijs������2��/�<��2;s8�&��	&ٴ��Pl�a� ,����6�5�k��w!��'jZ__��M��ME?u&;�@����0�!���U�`�G����\SE8�Y6�'�-9 wDs���C�����䴮�_���W�ю�\��t�*N�;]O��Ru.���2�Wk�3��\��������e$�t�N�x�c�����d!m~���^�c\�ʗ�w�6�5z�f��S�I�g��E}��1��1�`#������玒6E��3��\?����-ՙ�:�w~~����j�l{iqi�_h�����@�yC�Eoz'�(�@<fU����{ҳ�ot�o�p��������M#M��ne��|Al���$�Q�j�@6'8ѓ���L�_�.�{������ŗ)L3�q@Z	~�=!ζt?(�x~9vGk~<�6���5��Uf�7�5O
�}T>�h�_�[�w��&:Ws�Ж���z$7u_��E�@�v"!p��O�uyy��}��/b��|6���}�>������	!/�1�K?#�`��O�>��o��lm<������McK��e
i�I�7��Z�Y��Z�:�¨�?v��2��s�E���	ٔ>������P����������F%h.E��/��<���+��}�/���84\Ĝ昛A�}�"}�-e�)dc���u�s`_���c�%	��lQǲ���,�W��=�{�0��&a����l��Fce�Y��;�L��u���5C0����}fQ�n@Լo�8f���:����=^u?84�̦*3r�O9cJ[��D������9�lA�U�6�<��%놮��_j�\U�h)���ͷ ϼ�c����r-5 ' �6M��M|��m���ƭ�3�W��#���� Ǥ��Y�JT���'W^m����������p ی#�����~�E?�׹E,B|k���Rc)�t����`�2cDiv�8�9f�F���P �Yn�~�h�/��c�#[i$�y/��B���3丰4+���t_,{�^q��ś��8���F$��CS�� x��F�բPo��ذ/��E���U��	J 5:�sf���fX.v(��e�qo?H��`��=07m�p@R�������E�J����. \ycB�G�^����m�$I@���M�"��J�Mh�S�d��u�Ă��wڵA{�;lr�C�G<���dV�8��>��t�q��Zi���?�mEno��`cR���D��b"�������MfKi�{�1�o9�P�H���4��G�47�������R}g�F��hl빮�	oWb����l�W��
��X���L/h=�)��ꫨ^��
�"��I�QwE��e���r��F2��rEtŤ둾�5q�S����꣎�ƿ�}6���Dzuǃ����/��0 _E��~�I����i���g�@��f��{0�Ҧq{9�ɚ(�ԋ��WX�t�Q�]���	ʄ�j���ߥ���\������5=��)����3M�֪ۺ�oL{^P��eN5g5�'S@MJ���'�l� ,T�S4Z���< 5�)�8��K���6ӂ�m�l����S����O��'m�h���VT��;EJ�v#��j����N�Gέթ�����bh�������@�P2k�w�{q���d>ϘB�2����>��L��l�k�f�_W��?1[�� ��*���!����ɳ�5H�U%�qK��6�H��غ'p�|ס.�!�.ɿ�Y��n�f����I2�$�����)�1v�=$u�>����}n��`�Rj���C8\��<y�q�>�Y\:�3*����w����AE�on+q���V�����J8���A;r�50����5��Gt��)�4q�>E6�\����Ug�>
�Ց�Lm���N 5(_���d4�+Oh_}9�@Kz��u+SJ���]m#oj��������s/^ �k�q_6�&&�L@�� X�����?QZz�wa�ʄO#(UJh+��t��W ���(acv8z�� ��� ��`�=.+--t���O8��J�������"�sI��.T@.3!q�NQ +�$����3���Lk�%2��9���(�kz֠JT�9�WZ6ү�=H급C��	��ɬh��%�dظNi���5ީ�2E� 	`���v�Æg�2�F��U�0��ƃK1�a	!@=�nS!V���Y�Y��d}V	�\d�=Ga��ɐia�U���7�fD��VgK�lҊ����zW��y��x��1c}�48�� }.i眑U~r�7���+'���܁z��� ���?]_�f�X ����������'�{  ��(��nd�w"��8�{���?�"�/R4���x'�:P��t� �X�w��/lUl���ְd��~1#[y�w&Ɍ��dDk�e4���H���Y��5�L�[���:̆�]�d&�h���SM�Ȭ
����boOY���".��Π :����v�avIs���.z�\^��3�w��)uTm�fX���|*
���9��Ci�>��a��z�|�b��w��A`���&�|8���U�z�ߦ�u��p����5Z�$�0IV�Z0����=z!���͙̕����I�-�O��G:�J�#n�Y���)f�e�}�!�n�P��G���w��������2<DL|)(Ee6$���>CTMX�����6������$^`��8#���D�� %Y�7Pf��xf�zm�U>C��IՊ�1
�4] �������M�
�C��(1�G�;Q��8����U�T�����	�L�$�E5��*�yNme��0�4س��^�q�RR5�P]Y��q'>��q���ڟ['Ȑ]>������=���DhY�<�Nd*MÑq�����H;�&�஡����y�����}���DCip��e���W6恅2�����d�s�x�8E��ͿQ���E��\2)��Ρ����P�%l��Z�u�CiJ,�FAv��[�ye���=��-���V�z*��w�������\.�%�K�N)j�m�I'���+��E�����A^]��A�fŎ�1��Έ��d���"qeH~�*�(��yR�+�˕G�+�#���,��I+*ߨϧ�A|��2���%��6��۔�xѰ�
KY��F� ?6�i^䨇B�ه�^jd��z���Y:�X�{����~1ŏCO`z���`���9��=4�9����z1V$TB%V�k�!��j�r2Oi�z0wկ;�!ױRVG���-��H�t�Y�B�;��k��!ĽDh�2�r54��k����Β��M���S�ݫ�%pk� X��©&#����ǒ�0�D´߈�A�^8P�W�PF���*ID�i�y'����qY	9��7�2e�vEZ1e0+��(@Up��@���v��Fq_D�dH��F�y܍K�YJ<	s��vЋe��L�V�J�ht����ܬC
/=3��qlErn}��]��='�� H6b?�0c[�m�� �)���� "���F|�l#��3�*cg֑��|����Q��Ep�#T�l��*�p�����p��z?�� ��`��gxv^�1l����/�Cy~`����*�(�<$AI�(h		�$oOή�?'߃��� $E�w��ӿʹ����N:�$���H�-�Fj�
/�[����w=P� �u&`i?J��d�aݽ��`"g�ޘ���v���$�c�&\E��C����Vi�n�7��i�G"�ǖ�:�L�&���6�od�L �д:��/��f5{��&�=���o(�n����~]�V�+t"���2	�.�|>��{[�ԏ_Y�E��0!�H�fn�s�>&��F��iyU���X�e�eJ0�(K�=4�w�����<vI�M�ւu�do}+-dV��ԛw��F��ȫfۥ�2��/��eX`�:Nc�X��������_m⾫9~paַ�˜��v%�2`����[��7�UքR��'�MN�ˬz!��J�3C�D�x��p�����IHX
XG�ߒ�$�}�6Rmu�-�k-~����Ui��Z������u��B�Ŧ��:)�O	s����Y���ͣbam%mJ���\��Arׇ���m#J�B���B��߄��n�2�a��!O�X,��uݦu�{<�x�?�QK-A�wۂk����o�5mk[�V@���i�A�@�Q+���Z�v+7��x'�1�%�b����nV�	~�%��g�nn]�F��)��*&<��CyYrX0��x�] ��[m*ekT��`�v��=�uQ���1LD-9�j��Dp��<��i�|O#�_6�:���I�$�2��?�����&r^d�������aU�Y�7;��l�f�g57��y�!����Q�����'@�r�p�-�H��fQ��N>+,3ż&��#5{❗�����+���}��Z�����������3��K�%U)�+��{���v�����&�_�gb���8y8�sT�����S�c^Z�˕�7���+yc�b��Ո��B�0�Sk_�S(�{�h��-�5(Mg���/�nkA����DYo	� �-��V�hBW��
J�NN���38� �BP��=Ye����4g̛�(��uSib�m��u{)�k���&2��?˘�+@�e��k�Eydmui�5��{��D0u1���i���E�R;��N��.~�,�`Μ�x���[�>�#�*��#�*v�	�?���[J��/���+.�"�4+*�➺�����HƂ�i�f�yN���ޏ�%���hm�(T�c��c��i��� ��	�n �'����X<����	��O�?�@�[x��4��7���p_���zq�>&�Y�}(���6��n\��@�+���rHW�/�E�[w��'���	i~2@PĤ����^w�[�$����|'Y�Q�nðB��#�n�I�79*��o�%�YuX�y���O�����B�M���knIs%	���7�/
�j�|،�޾�c�U���J��D���g�ڊ��ʽ�+-f&p�p�ȅ�P=j�v
���Ľ�A��b�<-���ř���S��ʞ�a�k.6�嵈��>�
���(J�QVAT��i$��f��F�l24�h���vd}�2O.@Y�Ə-�A	FZ2i��nCNQ�֋�qC�Q��wԣON� ����Di���lS9��d(�(�)/����A�׋F��g�L�O��_�O)�1굘@Q*�B�P��ȿ����V������[;,��
"|M���H�l�M��d/�8�]-7�n�N��"4b#�(�]	TUu��vj,(]3hy��6Ӝ�58����@�xY~��nC^���m)-�gF?Cv���1F�_)}��2�z�D�t�2�${&)>'~��ĵ�q�*�9!UƷ�	�tN�C8!pԵ��f)���"	Q�yW�6��(J�T5�&�lǬ�wlp@UOm�2�ɕ/�G�MN��U�\���C�P*p97�@�c�I�|[R�vf�C�.�oU(|�#޴�qv��g��oא_� fg��PV'������ԁ��C�~C|1Y)g l���'Ӊ�����Č���|�L�(ֲ�vo��~r|eS�0R.2R�Z�B�?iS q1�1��}�� �j���ݫrz�?V�u���+.�b�����>-њ�RMz*S�
�o_,�jL�.�L��'-(O�}#�>Γ��
\�r��IE�r�����1n������:�owJZ���r����[�h��:K/�����(�"^;�O��f8k�6_ٻ�<��E/s���SB�� @9bq+�H%�LǙ���_�PBk-�?
��F���Qn����$�2p2Gyء
/>��x���{������'��܅�nD}�wJp��@�qk+=�3�d8^�cQ9�ġ@"Ə�Ƀ,����
��,����14�x�h���zˆ�	F7Jв?��j�w������Ƒ�t-��L�o��ͦ[�Mǋ�4v��7���6`��I�iE��3�\{�|����m��v�Ok3ㆇ{��s��vuW��J~R�)Y�0C~��KM����~�J¸���`�����˯s"U�P���L(k��=��.���7Ȝ(7X�����J���HNZ�܏� ӑ �ܜ�X+���.�x+���9`��y��"�y{W�`�,����6m"TE�G�H�yA�Bta Z��d��c��!h[��E.�O��ķ���i�7���]����q��YC��AW�Z	 ����Ѫ�U%�N"ܘ�K�%����0���F�F�&y�ݾ��+�L^��
�/3�yT����y�?S��>�CZ��߫Hj�X�w~�e� EG��x���m�,��86��8Z$J�[*�Pa�~i�O��wu��_����ߨ k�Ď�\P�Vݗ3�H@I�����$����s�t���54cܢ�G���0Ft�,Òp
�����Q�#�����H��ۄۑ>\����V�`��T��a~X�y�r��,���]�ã��U���>�;��t�ӿ1T>P�c�N������oɒ**ronLK���� �&k�c��2G"�Ζ�0o�A��$����~`A%S�����ܼ�U��:?.-�-G�x�?�8a�"54Auȹ?W��@�foX������ C/�����8f�>:o=y��u������n�.(.gb԰�� O����C�E����`��!�쐺��9�f��*��(�J��b��R�Y�;>cp��Ŏ��R��W��U�Y��ѝ`oyS�O��=�Ul�oy��g.	vP;���?!r��n���f�'��:�	�
���K���a֠^�hA�����?�t�.�%��K$%�^��`Z�3��1���
��õ*FB2�*����up���#z�hm��}�=J,�S��;l$���ջ�
ǀ,�=��r����Ԡjo%�*ɇ�������P
Z1��#�S���ۇ�}����>�t��z��F����̙� &�ː���*'A7=`�sޖ�{�	Y+�-Pܤ�8������|��a�`�@� !4<�M�� ��^�:�l�Q���|�ѕ{kh8�/�������2y�FL�T��r���^��gp�"��	����D���vX�qBh�[�i��EF�D ��W?W`������.ݒ�
-Q��"|��Ӄ1�ځ׃l��>۫�p1�1jNf;w�W�$�kWN�j�ɧ�w:��8����z��P�9�z��H��h�u�ч�-�c[n:#�m+�M�L�u��zn�����yh�7��l�;�������af�Z"�3(/��)�V����j�֗|s�^�f��2�s�Ò/��.���@��~�˞��yK£`ě���1��dD�gј5�j�f�R���x��6��R���&�m��z���[��<<i~��/jD���\G���9�5�4��5���#�Ư�Dg��ߤl��;u&�|DϚz�i"�����k>��&��$C�L��ͷxֱ�p^r���a�U@�.�?LJ�>�=������?
��2��õh_Q��rܻ��ڿ<{�N�<��\!'�Z�$��t�y�3 �T�	�P3!L��bm���hs�L��@;�
���eۜiɖj̬u�MZ�d��~�Ӎr�HW�΍�6+-�seA[#�$Kҿ��`����_�(!V L�uP��A�J�?�s�⧣�W��M*����5�y_��or�[���/��{ԐT��G{�o�wP��+���/�:���j�����i�ܛ�W�P�j?/�x��ѭ�������8xҞsM�a=��7M��@�
�Gp��<��(٨��\���]�s�΂u������=�J����!^us�w�y�#�-�}�~s�B\FJ�)(���	f��Tx@ső_ݾ;"�� !�S4R��g�8*&�/�p��;�]����H�i�3����|(����t��I �|a��+�"%$$�P0ザ�y��8?2Rm<Ĩ)��9�V���G�KGYx�:�qԧۦz؂�B���=�C��r�ԝf�q�l���h5S�f�m�EU��q1��\Hb��bE�$�Ds��� ��,I��G1갏��({.'� �L�~� ��`�5!j�)"�5�r��?�����xe��24t˱��9,bA����:�ϱ��X�������Ɍ��*���B�v!B�!�_��O)�Ǎf���]����I���&�6�H�ׁk)zI����:�#z��"Mf����{tOg3Z��L�E��0?\�g,����DQF�v��FH��w�A'�<L�\���X|��w7�e�1k�z�m+�D�a˳f�����\q�>j�ux<�n����6>꓌���n�ǲ2�B��x��}��05ط�l|�!<�	m�x>=��x�;����VP��un��_ki�����+[*�D[)�ں�q��+���h�r ����%��8�K-��	�.��kո��MR�nxw[F*�!'��tB��mr
�e"�A�>�)�'�/����J-�uD��̱Ç��r�ޞ��^'�c�J��������U��F���5%9�^����H[߅����r�.A�p�w��������G�e�?R��}�4�NG-����M���K����("��g[ ��=���*u���z˥��	�0���B@�3%b��(sڄ��b����^-�m�R�4�

P�6���Y����dd�� �sh�4�V6!X�:܋S����3��R&!�)6O!��tO�u	{���Z����8�l(d�Y(Af}/Tʈb���c\`.b;S����㱕9���L�-!���;��Ӽ�����2$˼��]�q����?@����UR~-�)�-֝����\]��y(d.�c5e@����{`�\���	����	N��5�_�a��/��v��E	�}nC��G(^�u�3$[��4��PH�@cF8M	�kW�L�%)ȸ�s�E��Xl3��RN�|3�Y0z2��/��������t>�};���+I{��#�lbOX�eD\/���14�h̖�+X=������C�v,O��v{�&�2C�*���^��Ս�L>�����M슴V���3"�=a.�p�I:RW�*�m_����n!%�On�<F��߷Ҍx���i[1G9?��k@0rA�P:՞���� ���%�AfVGUA���A�ˠ�-�oڒ�@���ŀF��p���;���9c�v�C��2�8�,�B�E�Y��7xBs������F�����_=7!o
�un)q'0�J"�Ǚa.���)Ԃ��ڭu6���5�oh��5/%l�I���s��֫,p���8#��񌈓|Ν��"}H#����|>X�B[CaU@���6_��D���e>Hb�^�(�R�7@�id���A-���^���U��y�G�$�_	���Ĉ�)�~'C
�W2%d}!��:OTyCvΛ�N�
z �_��뒞�g7G��̘�}&fM�+�2S&i�S�1܎ޣI��',D�E����T==������NG.�c�(�f+q�٠�c��9{��N"��NM�?Yi"p�H�!�6����&��]�Wt%�����0�ͧ�,����!8`��e�f�#Bz������I�C��	��g-�k�Jr(!�?���Y*\?�v��;E��Y`Ӭ<},O�Y�z��{�99���nup ��.�m5-g^���·�� ��n�v�?@uYZO0��ǚ3��7jR��6�ʃ�R�1�D����!�cF�۳BKa�7ߋ��R���.�v�K�^k�J�M�q��+m���_�(�2a�M�P��S_��0"bP���B�J�X�v4��FZJ0�V������솷�Hïf��O�W(/�MI�P�\�]�q?@`�̮p	�� #��8y��I���׎�%���CӚ�� �zQ�-$����֍�bc�`��WZs2�a;�0��T2|��VxW���jXS�� �#�t�Tܧ��K�@�$vb�x(�� ��v���	0��qf{7LL�~RsmP�c�J>�����ùqT�/!
&��ʐL}̦�6��I?P���l�<�{�6�B�`��ԑ���"�V��3���;_rn�����Ec�>;��c8�)�� ���A�m&V�,(��)��g�p;��2��  ��t6��̈́�Ļ?,(8�|Ԡ/��k�x
�I��~��$p\���"Ǹ�!�m�������+~4G�/F�$�H47�������E.��d;Ľ��j��xw������m�f ��<w?�V��[�()��M~S�#+���h-F�$+����� S�|�C��4�=�D{�eb�%bM�v~�(4[k2~P�G���sl��9���0�6%�%6c-mr#�x��@�&��c_e��l�z���]@k	�:%6��4�D��?�-\�����ٕ���o6�:`'9ʥ�=Z�C��n_�VS����F�؄���z���";*"��\$L~�qw�}q�ξhie�YMK�ָi�����"�;�����'���@�*��D
�n�K�h�08Ff-c4rH��k����l��G��p�Ɠ���4�2SlYH��5�3W�p��?��hh@B`|8�k:��۫�r��dy0'�MxzP���v�GՕj�?{�b�%?o	��G�G����̜��cE� ͙h��H�'�һ�j���&w<�|O$���X��\��+�'{�`,�6��G�4��3y�W���!n�Ղc�m�ǡ+U���q�lN�W+牋e"9+`��ڔ�)��h��?��&�n����1w���* ���$�ۛ�W���Y��oVm�9g�k��Q۶��Fe�lܹ҆��}
��R�q�_&B�&��&jm�P��+�<B(��y�tSA�{g�o�~����Va�-Î�>����U��k5�G)����l�w�h'�A�� �_���o��rtV��#�� \�S�M�T�h�-�Q�^���9> �Z����˶m5h3xX(ģ#�f�a�°U.�k�2�j�4���<J�&�X�TEMJA�����bG˃�>��h)�_��u� �=�Ƿ����ꦹM���gR$[�4O0�36�2�"�@���Ex(����U��'�_��I�=ZIM��rЕ0H����K�V-��Õ		�|�fv�ä���c�}V���\�V-��P�����A����*PRI��`�e6�e;Y�[@���ݧ��5����4�&�9����~[�����CLɱ.	��`�}3^��|�];�}�QO}�_z&;fuO�T���ߪԮE��\2��ʵr�ʧl;�I����x� �N�m���O�2V�i�����b���B���v%��A��؀���/��j�oL�X�N尔uP�́r��M$��^��o���	
���H�EF�t@m��3��PF[��;n��ݧ<�>	���m�WP2���-��d�`[�j����Hx(ه��S���]#v�gs�8*0@@�_�fk��8Y�c�hn']6Z@h8�WH������DՊB%�"��=�&�����Y���0-�qzSj�m�품�2s�tT�&��b��z�V.���Iy$�jTf��GZ9,�F�`��\�Cjp+r�*J�����dP[�.��"x�P���!���ױ��l½u��i#���ݱ�S1�OoJGч�� '��"�n����g4>{s/�$��]͖A��;T���+7�뢍��3%7����)�e�W#.J+�BL�&c�z�U�ۥEr�������m7k�\���z�l��A�H��
��ދ�|���	�� ^i��:�G}�zn�M���]��[���:��?��C���_9��V�n1WeO7���I��Zʬn�"Z�P�����]�6>=��LIvr���wv�i,+�&.C)�E�z�o��a E�&i�^�2� ��xé�{U4؞U�h��ȔA}^	Y��5�G��O�y�����/��ȩטW�mF�_"���pf:h�%*��A�|A�fƓ-;#��UpW�Sl����? �a߼�{ڶ���֎�>�#~��a2�os��g��z�m���{#K\ǘ
8���a������UDG<�n,�9��/S�`�[��{.a��lB���V?���Ǐ<���˸���z���M\x���N}�?�Lj�أ�('��n4�����e�h��š�@�J6l��W�R_/Ri4`X� X�\0���a����J	,(��a�d�w�S>��b�(�e��_�-��η�����[j��<�����j2�}�9�:�L�ULf�YsW��������� MȻn�KIe�~Ei��k��Ă#��8L���<�t:3��Ǐ�W��9�I�H�2h�Qea� ,B����cd�/�8��t�0�9��o|���A7�FaU��'��^�W���<h�"�iFM����J~Ɠ^��Խ��?0��I�^U�{B���ǒ,5_~Y �KUl"�L�S�l[��R(�g�ſ@�%��-*�p�gӚ����L1x>����H
߆Ar���{��Ý��hEJ7O�Kx�~�Q�7�n���FE�Ȗ
T��b!�
�������m�4�'�%�r���N�<�� �`�@d�$n�L�t���9%�h������9�=#\�B�����je�"H�)���o���~=�ٺ�G�ϒ�KEʶ���W�nlȒ��$��D�ę� � aW�{���6��J�?���p0���/�&?�B�	�n���y�P��[)�Y�N�� @����"���P��C�]�ò����f���\b��3>��jQ�D�0Q� =�c����l�1o�1��\���7�2j�+z��_�9Ђ��[�c5%��z���A��n'�QL�*t��hp�����ߟI���h�e�cb.������%#+ ض��"%j�/��
~�RѬ�s`6=T\,W�D"I!T�9bW�ը�J�?瓒�b䖛�_���bl��l����k|���R]�xHsU��j���,U4x���!&�RI��,r@I����C�m��cps�Ѡ�[�/�P�"��{������.?.�e�5uN���2@��_�HvL^�1�&š�#���?\��z8g�z���I5urT��o%��E��-'=�nx)��j�	����L��a��3A�gz���i�K���i���+ ���ߥD�p���7�� �
߶Y�Zg):^�oIX�aڢB��G�2���9��A;Ȏ+�J�]�vh�튃մ��]�-`z�,]�$�?��:�κ���/�V]�	B�Wu�<�_�]���{��L?�I�ԈfY�ޢ%�1k!�a�"���X��Y�����"�9�W�����y'��V!Q�s&{��YP�W��
���,�L�W��/��~?���!f��2$���z�瓾���~�NĠ�b��QIUt[�r���_p��2#�rB�Z�SdnG�5 \��vp?�暻i�m�!��|�͌���&�z'5x�,��2���E����vB�^bM�B̤yA�G��
�{��q��,sߡz��H�ƸR��`���D�+a��Y�|���-�/9� �ʖ3�yD���_�A)M�����+_ۮ��z"bi^ ������'�ߙEC}Rgc��v乊ʺ�"��V�99	��=ָ\��K!5ұ2�Ѭ��z@l�^ݥ���9%T=�"�l��۠Ӊ���pϟk�"�C�Z3��f���IH;�a�9�iit�)�W�yg��ŀK���x����?FQ��fÍ�\��倆[J軺�tעӮ���v��9�8������v7(�[ָŋ�1�߹}Ϸ��m���xh���䈨x�1vL��{
��b�"r�(���U��%��,�j6*fk1�m���([�$��<g��[ZZ;JW�Ӥƻ%�?�~�þf&�{�$�Fϱ�W�]}vR"д\�� ����_MC�CO���s�x�쾚��-C��n�X��Mj�9z��k���(�0�XC���f�҇���Z���$.ݱ=�c�a\��2$�D�`�j��r��w�?��D�P�U|��se��/�3�15˓�z�ڰ~Y����=_U�A3�>OL��%U?�W٫�]çi@��W
��'i��P��B��Rw=ޒ����m�.����'�_�aq? ��V��ĝ�B��0�I!F�x��-k�NXD0nb�Ā7?�Ui�|C�nȰ�����=CiX)+
�M�>�Ҫ3�X�.]�d�^1A'�T��n�42
�b����{���r��D�������w	zO�Q�ad��y]��97����^:�z�,�� �K�e���Z�5-xFw�XK�D��Ha����lj�*
��r�"4��鮈�I@O)a�aT�o��tB`h$�݈�Ę����'z 89
�U#�=��lf�d�7��3k���׼[���s�=�<�v��յ9m������8�����;l��9y<��J�����g�0���_!��z+Q�{�o��evmR�6p�3�cN���2d� 4}��Hy}�ņ+qU:ˍ �-f�B��t�G�㾛dפ)-�{�W�����s��$�U��q
����-ڲh'��H&�ϔ�
o/�.�`��(p�%V�瞼��w?�������N����4t	�#SՄ��J���v���%WD���nF��jp2.���l��,[�@�P��\�T�Y./�b���Z�D�ueA^R��i�vf *�M^'��w�9��$���˰8R���!��O�Fa|}]���lg?Sd���\]�Mc��Ѭ����$3m���q�K޷��:c�Y ��i�ԛ�;�����ˏ3�nH�q# ����W�88Ų�f�<�T=6�M/O����m��ڽ���������<�6){q�w�r>
�X��?�B/��1qǐ�+T
0~�r.J�����V݋�A�M��P�B��
W���T�2��e���E���L�iB��x��\����8������xST-\n�}�i���-�q����]�hQ����3�F���m߽GN��W����������d6��o�}U�]k�3P\nx�77�b�O�������XCRtC#k�}��َٗK���N������,а��O��\�����"ѳ�\���
��Í���щ3� [�0���싘�E	h&��}i3�!��ʿ�����#ԑH o������
��(,��ъ���t;ak�k�nx���I�(�����F���ص��%��]�3���,�]AE���'8ZX
��M< �C�ؖ���cg�,�R��a� ��7��=����X]	�]��l�i��٩�����R�$���=�D����D�eXYt�*:v�aOi��T"���ш�{a��l�?�&J��
\D�(�d,%��\����=6�����iY]7��g����fC y>�V�$�j7���&�^z *g���$�ހ���i��#CϓE�qQz1[_�Õ �3�tP�i.hk�����Q�>d����z��S��6EͿ��YؐGPJ0�c�w'ϱ�,�x���%i�Ƙ%�5
]��Aߙ�@1��,@R�ݣ�֬�6~cGB�cYO��5�
yn� ��}v���Ǘ��5�I~�o��z�	�-鷾X���'�E㣂B�JUz�n��.5�q96mI�ט�c�pu��Z���,c�M+n�$����-z����6�K�|>���;k���>_������/:���<��]�x@p<Y,~�]����c���:�َ�v.��焸���{�[��4B�w��a0`ne�Ϙ]�ى`�e=��و�ѻ��D��m��,NLB{��zEP�4����;Ĝ�"d�tW;��j�R�B�x�._8�t#+�%��l��A	�bG{x#��&w�����EO�P�h�Ғ���[5%��[��K�$�gsJQr�:����6�#$^���`�]�n��UO�W|�I�����͒�u;�;�\\�*�wTWV�[2�~m���U�E�� _����F�Z�-��;Ud�(|��上*�bRR��#�N�� ϻ�pm��ݏ���Mi��K��Z�s]%�k_���,�%C%	3��f�.��1�Z=��:�KE�@�FC��0��L��UHֲ�4���cA���bٻ������|*����_�>	O5Iƚ`ޝ�d�	:R�\�7e�$��!\����(�'H�?eOI���ٮ�	��c��=�����K�Yfh,6H�Hwׂ ���F7"�QƩ�ݶ�5���H�*rv>ꂐY?|�����7���kJP�M�����$��pg�=��y��cpv(���ٵ�mG����U��\�ͅ;!�	-�JC��̾ӗt&�\��<�j��|琒� ���ޕ���я%��%�n^���Ҭj[^��x�!,�iFo��W1�Ud�G�^�D����������Ȟ~kɑQR�uN�Jf�!��]p:;P��܉����pO���'޽"�J��4������C��֠��"��[�|U�p�3B4��-c�`N�<��8t�}$�����q�%�A�;<ݵ����v�h��;;a�&{c���R�r> G��{���z�rN�lX)����\Y,b�Q27K��!X�P4�5[tW]ѳg�Κ��~j!����lfa�'!2'�qm 2�рjJ��O��@rp��a�ft���u�����q��@�i ��a$���S��w"YNC�m�Ì�l�bV�ƕ2����(p!����Yz��^�T��Qj��-�B���ٮ��a%kmLSO�Le^�<6;�B��˛���\�����t���6�%n��z�I�^c&ʖ_p;0?���kb�ǨjM�ee㘊79 ��:	��(�ن��56ѥ��l1�Bp�6h!�3�DkI�H&Z�G�E�th�I%3��<�89�6;/�A>:�ԧ�Igf����Vc<�Á�+-ʟ�.R|x����C��{+��zq{̐h���pa|@K����������;�����f���w�8/z_��ʌbH�ӣ�"?��]�^DԔ�ᮋ �MK�1��U���EN���������#@�g�Rz:C�kq����m�\@Ĉ��G3&���m 77~�/C(�˅�Y@��)����-�<-W���u�N�]R�t����`���tX��+w<�:X[$�=����MN��0E��^^P�҂��bʃ)��K��]��Gf����D��aXxV
��m�7f)LNY�;
�o\��Ԝ�"<B�T�핯��gV��uR`������/��CRѪ�G�n��c׳�.̽KCh�u�|�_.	�K��$�,:'�flf~�G~]�l[�������j Ȧ8��n�'O�����g��ė =:���������C�K��҄.�����ܱ�3ix�m\s g�qR��4r�x0\�;I�ɖ�Co��;
?�~��H���A�u#.���V�*�J;�~�Ľ��?8�r��ܥ&�T�7�@�nC�ro¦xK`��o��T\a.�_r�pE���jO�C(�� k93V����tk7w��)���H_���iYm���w��H���:�É3�xᄰ�+�f] �ԕ��LK�Yu�l�K%
�Fѽo�
��V[h�����E�a�6�����ŧ7�q��؞�Y��SB`�j���˃=|���O'������
��U<���FmԿB=$�4�<�۷ѹ��!i'�/2Y�����$��?}=;ʗ����yOV��3/*���{0dD�9@��o,�2�^ܺ�QboDfgl�� ��GG�J�&Y.$m�i�{1�����FG*JA��X��p�7et�]�7Š�إ�hzHo!�H��5��K��}?xa� ��e�	=�8��>�颖	�bSh�"oQ~�f�Q��D'�T��l`���w�g�he��C��GZ)�kTr�$����3�綠��\�k�l2�͔V��9��\�4�x*	ݔ�$5��
b�a_��$c��1�,��}��-�ou�m�#�vO\�Ԟzr�?�3��5���Wpo����O�Q">�2��=���}�?G�\<ncX<��H~�?���o"�T3�\Ljf->~B�D��}� ץI�RIT�Za��<4��&�ZA��8	����H<�[�c���~qI����\�n�&���ihiG+���_|M/���|�!�[��P� �˱MΖ�����*�3*[��ґ��N�d���!5J۸����$��S��;�٠�Vy��uxW������Wr�f/�yF�ݹ�A�_h����K��Y�;6�F�nЙ7Q��[1K���l���(�
6�O˔�/f�|�F�y��r0bc�v�"U���4N��;��	N����k�gfI|�4Q�꽅^�bE�Pk,Q	�C����]�����B!u(7���44]<]v4E8�яg���[0���G�uE/G7+p��n`Vp9�W�ڵ����S�۰�D�ፑ��4���N?[r+���KoZ�Lņ�[�$C?n������+5�l�w�ǹ7M|����{��;���K��z3�4���X�cb���5Y��%t���Wr2ˤ�-�Śړ.������N�l~�w×��X{2��ۄ��æ�$�+ �9�n����dyhaM�S��)����J�#�0��yG6��� ��3��B#�O�.��	+�qoĪ��Cp3�ّT=�(T�mD6�*O0��? E��:&@=	1��5��Ԅ*U�������G>���c���QM��{��y8FZ�gz��:pW�8֞�9����;Y�^���W&r��K6�"�Bp0BA �x�q�@�4:�VGSN�Ԕ<�1T����ѭ9�1��S�vk�s�F�n�&�2�&������:j!���:��j�Rs��Q	�ϲ�Z�v�iw���`FC��<�nM�i�U�5�������V�^kӔ�d����v	���ZXj��P��L���ՀWߩ�9fUX�n�K���$�@s{l��`��-BY�l��j�s�f:1�M��"������|t�W�f�\�6�$�k�YE,�C7������ �3�B���^����$�f�nN�y��i)%q�� ��)>����͊��$�i���m\�C�S/q�[n0���T'�J2���>Z��?<�jh��R�3f0�/+WmT��f���(����?�����WZ@�E9'yi�����f
������ݼ��y�\-�$���	�׹߰��N)�Y�D����rZa���N���� �*��5�S�"BJ�~�����Z��`Dɴǥ��ׂw����Φ��LM&�!g~���^RU5
Q�槠Ft�1�S�Gg��j�X9�٣�q�.WB�H�O��%�imc\��܂k�m��7K��q�/Qa�]	�f��5$�u��qLf�R�`��g ����$h��9��C��N���e!]��\=��X�I/R�5�8d9��p�do8o��D�
��\V�P�� �v
�E��skd9(^S�n���i�ã`2po�뼠)�M�tB���y<�������}���)�������f�M�J����N�	�#��gAf�*ug֐&��qTᄫ@_�)Q�^����:����"�#�g����c��u��Y�4��?�m� &%����Y�?�V
�������=$P��Sq�i+��������d���sHd~��!w��耬>�Tɨ������Q6uL@^��+�@� >��Y���5SD�������U��ܑ�(�Eq�H�=}��i���S���+Fa�*��$~K.悓�o/��L��K�_T�0�!�̪ؗ�ZB�lR���RoW��:����[*�V��J"iS�gC�2�e�t	�tK�:M����欂���ha9&����6�[�x�CI���C듕����ݔbH�`�_j��c��r�6j�$Sڞ
MAˑh�'��T~6VO�"�F���r@-����)���?F�I�r���yNa!��������&6�2��+����E�D�4���pnR���g��q ������j��ѽ�g2G�L�Ohj���^�h�LwbMS��XE��׺���q�.��Bc�D�Z��+���k���`�I�mU�C��=��2��64]��IU�9��"*������,_a��5,�]�;)���C%�΃ �0����
ƴ W��0]��F�_/�P�38(ǏxmL��a�E
��?��m���T��9\Ǘe
+K�N8g�R����� a�T���"��\��e]6|��H��ɱ�&�{�i\�^7��S�G#��݂�HSإ�w>�(��$��!���N��ʚ4�+-�F��Q�Y3��i�$/�Ww&\�Z�,�����U	��i[�ye��
�0�!���:4�P6����u{I9�P�P&+�Il�{��_�dH�Y�B�ձ�4N���%.����6i�]�V�ߐ��IYA�:H��_�ȕƈWF�;������R����"�qכ�@q���<B����b
�q�{9	�*�ȗw<�Y��c}�/l���w��%ӽ�Y���=y8�����Ų��X�bٞ��MՌߗ���Q	JQ4R�}�[�&Ϗ���E��$;��9�7/ߢH"���׸�yM�g8�]������ƥ*�	��j!�s��+�v���J���̷/:	���*a&-�{�A��� �{J�������]��
g!5������L/��FB���DA{́�ҡ�6�N,bϷrW��i��k�R�/n7���ʫ�2F���)4��٣�ep�=x���<|��8�2:�� u��P��v>��d�%��%�jj��W��U�F v?�U�[�3�[bj�rZA���;CߏJ���ph�i��кN�߆�����`F��+�@�ُY{�� ��J8N�|�JA x��2KG��Xg��������#�_��6μJ+�bÝ��G�=d��2�)��f����Pc�;R22N��6<�F�\���<��#�~-��
=!��+���7杆�cx�	-/�P���L�P�S�B�h_ы�Q�#�9�"Mo�������'�]�E���)/ԯ�%��۹�f�o�O�7�΀��2:���'y��?�c�:�e�X ��V�ll+�@�U�*b!͐�!0���3�@���7�$�/pG�t����Zwr\��у�;�C����z7J$�Y~�N�����T[�=E1u���_�#�)�ܨ�N�HLȗ�ԣw�,�6$�1,�4�����ɦ�`2�ݎ������#k�s9��?y�cƏ^����K���.E���M;[ ��G��TH����S�"j�ߓ;�XOH=�(�a�y [qp�� �������wU׆�=I�솰�%p����#ٛ�g=3N
���q�=�o[�Ձ$����o�4�q]�:�H��0b��:��w:AH~(�z��s-�0]�UL~Bp��[���w~�B��A������C�D����k^O���dU)@C����c�^�8�j��6�����Y�~ץ؃X+�}^�i!�J��^]�А�>�4?A�i�n�����Y7l*�oY��a�F�3����В�^8�XQ޲�|��Y��hw���C\��m#ذ�' ������l���è��aa�Y�8�#$P��ŏΘNKY	�f�`-�w㭓0Ɋ���$E�rI�&������Խ|�t,B�>cAR�ҹ�>=����O�ØZY�L8,A�=�~���}����Z1�b������f��I��Ge����&g�V��v�V	��o�k��!!���=o�$^���lܯeNY���f���ڸ����8M��˽�e|���S��*E�FѸ #	@����[�����@�+�;	t*�i<el���6�R�06߻9%�������=���]�� �)�/$�Ʉ9K��L��Y� X��k0��Nݍg���qF��h���Vm���5�%lpCul��X6cK����7�~)�'�ꡤ(�s�)��j7'���@��v��x�
Kn8������u�s:�Ș���b��i&�n�\�}���G��կ-n�~?�aCm3q�=S�#4�KIy?I��{��t�����g��2�a�"�B���Os\�(?}�N�W��!��q}�	�}�i��\���A>�+�5⮿q��B�p����Ǝ�`Fmza�X��Rz�
Ĥ�/��
��7�*��pU�>�C��D2��0����~�̇���e=��� �[��%�,Ǿ�y�b�t-Bt�_D��E�,�).;ؕS%�S;ń�K,گs�A)s��g���s��"��2�+�=��&�ӻJ0C�3m��x[�Է۶��<��j�/�c~A$�h��р���:���W�%{=��4	^�̱�g�ŵ��	��ƺ�� {�Ý��̵em{��r�2��g� ��(HNߘ�YWX�z�_T\���V^ۃﺢ���ĉ���+��-���?�����C'g=R%���̥U�fk��u\0o ��#K�4������������Q��n1k����?��R�.e`���(�σB�vEa��N>k#p�ݧdu�Zov��ǝ�I���ar����d�Kf	�@ኯ�~�E>9Y�������x^ء���J�T�j�.T��ϑ��l�>N2�5$�7���r*k[�N�N��X�����Q
KW\@I��u�/����������K��]��{��Oy9�i�9�,ǘA=���H�M~U�S�G�ɇΤ��0f��Pٿ5���!6Xr05G2$Dy&���U]<B#��;T��>���|�)�&�&�f��c�|�<���t��r��NL�2� �4�#h��p��^�͛b�B3�F�2k���Մ���A��np07堂��mu���4 q&����;[8��ɠx� V��4�Ѻ���%6@��4t�>Q���3� 2ׁ�z�)�a�A�ψa�Om��e�ΚÌj��틾�Ջ�j�&I�=n}n���%��k�r>����"ĵe�`�{�+� Y��PS�'��IO�$;r�U�0��\S)��>.��с���dg��h�X�Bu��>bS�Ow���h�P�i�kj�vtI����������y��& ��f����Q�h��
�C�b�b������O�H~Ò�5�h�>�*�5Uz�Vnѿt�>���\�zX�SX��v 1�"���>���|�׊�AؠW"���r��c�O��egx>�Ρ�.{m/��w?TT+�6��s�I	���7B*%�޴���;�@�Z{e���l/��ک�c�ѹ�>Z3�G��Jq�f���j�����8/&��r��1�zN3ը�;��hB1V)�y�ȫ��ڪL�4#�?�r�x��[��PV�}$o�U܍�Lؒ�<{��'7�;�%6��pɰ�����E*�L�8ۆ��"
���:
=pZ��$2{4]r7T�	�T�R7��F�+i�5=��ܻ�Tf���d�����K�.�EV�~[����V��
t�+��>�����GNf��M�_ʛ�J�J�~��k��/9�@;���VL[�x���da�0w�mr��
$��G%`G���{�#���߽P�o�!�J�=	3�ˇKmȡ�>���Sr�� �]�)ƭ�X{D�Qݾ��S>=��-�$�$eP����+#�����P�ĸ�n�>�[�$��?6Y'��UFzz��o��e�X�1_���S\�Ri�O#�� Қ9,�R�ߪ�M�E��B�������i	H�Q�Qq�z"e���O�NU	7�[�h�B�Kt�ҿ,:����J�p#���*4��[�F�`��aF&�&Oo`p�;h��f��j!��Z����DU�
���Kp���w;qӼz.�s��=竜�7G|��������*P9 2l)>��Mw֭�4�*��`���z�t�u��̗�;�y�=����5N�����^+ ���k�����Lm��WZ�*���r��e_|�
=����dG��ݠitR��B�ʎ۴6k|G��v�uY!�k�=A��j�N����0Tb�BfI���]r6�(KY(�v��cF=wb��;�uw�'Ǥqy�97���wv��?yԸI�5�TZ?�^��*��t�{�tY_�-V(P�Ñ�&?�+�=�e��P��y�D���0��~�.NH+MJ������5�I!d}Z�U��Ы�w�1����ag��瘽~	X���Q@(Wtf���,8 d�P�X�� �ɞo)m?�s�U���r��!ӧu�¦ ٜ��˽����<���-֛�cO1f�G\�i ��1�&GEn��3VV4#	N6+'�1���Z��04�#l P��y $�碘�(��xW��S?1�=r���͌'��9�~������	�{�u^53l���3��O�fQ���/M��g�_}�@���1��B���t���I���ieI���*f/Z�	�[�s�C�9��/����̦ל�'�Q���c�
�oqF��t�D@M���]�'��������(��k���h�j:�;� ���=L ����~�b�~�D��9��hAk<��^2�Kg��o�*�-NY�eIƚ�4���Fʝk���Ƶ+N�M35G,'k��H
����u�6ǯ���w�n�g��N�!���i���Ñ�pǭ�K���.pSR��a+eb�8}Z� ��O�T�y�t�l�p��2��ެ��.����CV��N��i��
�i�U�o|5���ܠ8���}�0����������/.�e��g�^G�<Ɵ�?��3�����@�؍��t�)��*K�`/���K3L���ܚ��@�:}�'�����a�dyl7.S�����%��D�����dD��� �9�*�U	��z��O�C��Ú��*�o�if	#�ݑw�N8�b<e�\�oɤ��~u�Uk�>=�F��B �ͻԅ�E��Ȃ�@�&6�o���pbD����Wj2�@q@��?����c�ʠ�5	{l:���f�/ؘD�!1�D�`��Sl*Q�W�Z�C ��!0�D?�Y]��{���*�4��0�#�#@I����iI=&њUt�z�Ei	_oSD����Ԥ;T�iL>��G3�_t�������6��e��Z���*z&�P(K�t'H`cW:���d�n�χz3r_MZqj5�D����K�����;~�h^����S�9�B���0�^,�d�_#Ya�\��D��1}�a� ��&P 1�E��3DK��c'V�,��a*��b�ނ!w����w�)+�P9��k�|�l=Ô�ht��cF���-��FF�8y� jY9����{S{��j���~�U����a����F���e��8�����-�n�9OJX�R������1�w���kF��:qI�q^_@���mm-&&|{��v��y�P�<PVև�+d�7j�
<Z�߻
�+ԁ��M��D�_�t0����B�q�
�ӕ��� ��]�5�R��G֔2��K�+�U�K$h�ԫ����ô���n�_�)�^/��4�=~�~�Ž���h�L�%�˜�l	��$(�#|Pi���A��A��͝��׼�s�LJx��*�7g����_y��Q�gFp]��ݯ:��7�͎�J��@�{�F���E�s(��h�d��ж�4�c��n��o*�%�9#�os�`��/_F4	4��	njE�/�u�d?E����l�����rT��4~:�^�Tq��Z��A����y��^؛%l�
Mh*5O��"_��X���Ԯ�p'�BkBu����� �vX#LcHm����Z�{������#�-�۾��<�I�;�L[e���M�_��JOi>�<�)�q�±i�t�$_�+o��1�k®B�U/PPdy��Ւ�9	D��}M���B(q�m�
1�R�<[F�ӟ2�^�۬�aX@��Oy̿�Kb;c?��)\ʴTd[C�MV��R�3�!�"��$jw��E���)GLs�֨ ߖ-;}5�V�A@�o�`RD�)m[Ԁ��Ȉ�aG�3�����"8*�ZI��z(�Y|�(G,����m�F��v��vsO�i�<e`���>���us���.u4�ƪ��d�y�χ���Ƴ3�c[<�����b�"Sw��ѵs����i���b�2��0�\�S/ۏ�'��B�aZ@qE������@~)�*���W :�Dd��jm5L���_�~�9O��" [�"W4��>W�'D�T�%�-	0����9�3Տ��G���[��7�������s� &��!<����N b��d#���`����&^�LE��j	���@N�lV�z��D����^��oe�_7�ʯ �v�� �^
�����W=�lbL���\
��N؂�{�ԣ�i�`)�n�=�{���K�SBO�ȷ���}�N[�����3�7�B�=�V�z��/s�좓�L@#�,�� ƽBs9i�;?���ҥ�ɚ:(�H�$�y8|?%E�{��I��B��a���~	t��T:GQd��?Xc<@7I��",!����h�����MQC�V����
����f�z_ZCZ�b��7쮙�ud�-�V���}�V�7@�Y�v zy-&������Pu�J������Ύ�=������?!a�0ҧ�F��w&wy���C������ S.CE�����{l����<�t%+�ZΎysJ_�+2&��8�r>*���w|^��u�=�Xi@�nɅ$ؤ^���&w��J��}�ݴ;�r�Sp��t�]5���潻��K�	�WiSV����+�r}U��[���`�~��|�y�\��^"����y]���.�5�H>������:�x�@��OH�[����jC�I�rJ7K�d)U(9*GpR9�1�Ȧ��!���x�w�s)��x�m�`�q�~�<�bC׃7�Qr��r��_��u

ћH�%3D�L�%70	��ۯ2(|����K����c@Pxt�ͲKw�=b���M��R�D%���W�.+�x�W�8�=*ʻ����W^�����UK)m~���Ï	�؋��|�6O���}��DPU�����bt��}��!
���C���Т��ZJ�˒x`Q�4DZ�]n8�'�}���q'�t��4�8���(�x6۟�5y��Y�9^ m�j1]�(Ҋ,� 3<�sΆ��Kr�^����߉�>�����n��?����D=Փ��ED0
�%�����$�'0�+9-�	 ʆ�+�
\�>�/]cX;HKL�2���]�%݄��L~u�u�"��+b՘+?��;7b������H�����>;,\XzI$��Kp�����_�չ E�Y
~�52��y,U@�CZ����l"|��!VS���#c�Ěr�Ǐ'v������:��A<�Z��+�[Ղi`Y���0k��f)��o�+[p$�z�ᴦ��Udi�(f.�F,<ɧ�^��c���=��!sjh�28�ۚ����b�t��p�+�X�I:��&T�����W�V�:��do�ێ����M;-f��U���M.�8)��8��]�Ԑ��B��AUB�+�/���%��$WȮ�j��ptH���7�%[��W�^�|�n@'�_-E
��{<;Z6��~��шQ��xU��[���{Nf>ۦm�2����P^0a�Mf�'C����}��w݈B������:hu�}nr�^�=Ca>�g� ���Z1���3�#�������-��{����^ק`
�C���9�sc,�2U�O�"��-xÇmHEa���GQ�eH�v�Yc�2�/��;(��������`��=7���^�]@k�V��eq��P��,3ݓ��R�����4+��h�A���F:�V�iS&�0F㏖2�6z�`���p��"Q�����a��=%�/E��������1�l)�X�0v���7��\,�y?pP� �J̸��æր짝T�Vo�<���i� ��b�������id�����8c��_�U��ݚ���ކ)���D�<��%<���zU*�_�q3)1�wi`3ř��z�X��f6� �ƽZhsUӗ"f�cxUb{|�:��;Ӻ9�O�:�6�R��� '��.nQ��X���+���&Ġ���� M�X�*Z�+-tl;��KWTx->�,�+N/�A����F���g�ߝ,{��z%����bL5�tȠ!���3�|�(N؟G^�8���5��?���ݢG{�JO�f5b��'(A�����)��T��$�o䩊�����Pl;x���G.�5֭�'z�|��m�;U-�<+����F7�,��tGP*������dg6��`Q0Z��>sMB�ԃ2-���ޢ6�{�Q/��N�-M�~.�&	uVN@+b���_P�����7�l�i ��[���?��8��)x-MA��r�Å�HL����7ut9��ð']�ݓB#�p�s.K��zj�Xh�[X����B����Ҟ��@(�p7��7`c�Ld�PV���_❎�D�p�7�۞?��읽�y�n$M�#:)�=U7@RN`U"e��-7�㓊���8��e���pE��-���f�8�����Ov
xE	R��rǿi��u�a!�'�� �K.��^C�Op�`S�ym����������h�_��� ��0������ �?&�@ Qd����`��B,��*��Rm�rG`�[�jz���J���}����1�'�)��,����fr{/Jo#{��ϙ�Ώ�L ��[�Q<�<~��y۲{˒��@�T75X����JEs��pY�+�B5p�\bҵ)��h�n��W��eBܻ��@ͳ:g=�z:�RY�C��}�S)�m�z&�$W�?`Ye
�ٛ���螀-���}�E���1���(�.�)��;JT���g�3��c��<#�t�3z!���W���臠.+���言5��DKt�4G����_ �bA[�!c��qE�$vEC{�ZǺڕ��d�Xy�(���jV
9�a�R�[�ĢS�j�4S����;��*�w��w�V��]d�p!�r��r2�>Y�����.#Ŗ���Y�{����e5s��|$�dZY���`D��	9����@gO�IvS?"�K��FS?�
���]U�Ӳ9�#?#p����B�P�[�06���$��W�NԴ	
��?�p5&����hЛ_�.�PFcNL��X"XM5�H�vR�qX��C[���,����q����tk޺g��s�,��,��jSԇ����O��C3�8���U���Z�W��+a�(�Y.��� w���SkB�X�-R$遺q��8m��ت�LVƒm�<�n��(��^�w�B@�_?yyS�zv*�&e�p��}���6��7m�ľY��˗8{�_�S����dTZ���gl9�4�����~G�J��q�~^�۾�Ԉ}�+�q�����͌r�*��"��G�*[��!àG���@��鍐P������7[����?k�($�\�4Ħ�4W�.T����F�s�Ձv-4Wn�-[L0�t��zN5��r�C���ͦ"~���� �X�Vب���X��:���{(���
��K�
r_�w�-O�D\�uQL,��iٍ����?_�uF ����H���
o5R�Uz�4��9���d-�N	p2�0�R7O�'_�7��C��KዲԠ�|�`��
2��óK|~���D�U�]t8�x������S�<���qN��y纀�N!Z��T��]G�sAt�� .�
�7(f�=�mc{tf�ek����Arr�"6�B��-������o~���|,�{�~�\�*���ႌ�Mf2���1U�IX��+����L.t����E,$�u�l��n�gJ�5��p���NV����唎Զ��d.t�2�s�	��)���J��7��L\~���6�n>?�#81�����CQtGK��Ī����ݾg�4���vs�V]�����.R_J���16S'	Z�%�y%s�ʷ$���u�'��Fr�Y�J�NK�o��"���@�*Ȗ0���s�����ܨ��P�3�f���L~�5 ��I��C8�4Q����2wӖj���7�ҷgR��_���ޑ���W'.ȕT�B�q�y�s����K��bޫp��xg��l��D`�
*���r37?U���:�Dܞݏ@w�x����$���ǳ���w�l�E��x�1Z���y=V�x ^s�1c],�7�r	� �[n�������A��H>��U�hH�d.{d1�U�
&L����<��q�F��*���/�|j��2��������l/.O���O�.�,�2���
)aTj'Kf��#��,a%�φ�D~�x�KH��qWn]��.e�:C�� �B�������%4����'GñW@����r:�ڜh7��S~�r:*<'��l	�"_ǩ��ٌ�8,6���_��yw��_�gc�%��[�/"�o2�t^i�u��n�ɂw-d�{)۽����˥�:�*f�V}JXrÜ��&����F~�=�T��v����`�j�n��7�iֆFS��^]]�Ī֊���y�F�-��I]g1�ﮦo_�M�G�N��T���ǻ��毒�n	x�a�&�~(��|;�/T�H1\͈�;��Є�x��D*zuc�7��a�'j��5�whn�N0rR*	��3�k�m��Pҗ���`3*e5��%�UnZnMN����N�" rV��&T6!ƈ=r�Wc0�{j��q�����l7��S����Bl�Y�1�㟄�����R�AK��ʴ>�+8���0`��ߜ�!p%�L�/$���0��t�_�e�	�����
P��բL͔b�WW{�w�Ig��k�xA{����(�խ4���=��9۠�q�7�nΈ>�JU�J1��!�W����ANk!��"��c�VQ��&!��~X��A�R��9b�_|�t:�*��m�y�T�ӵk5A|<,���(�W�hbF�dz���m��/$�Ԭ)$�-���<��`C����+)c��~��^��,y���<�������ԉ�F�Z��֪�ݬǻ��A�翲�]+J�2�3���Qz��:�G0e�S^5�S����P��+�(������	���|o`I�e׊̣ϯQk��1�S^�t�N�L0 �T37`���)�/4�F^�2m���x���EjP�<vZ�tvKw�]a�cʟ�a%�O
J�����������1s��٨�C$�I�J8H��R.'Pn��.����'v~�E*#�S	&�-׺M���-��u��b�J���5�������X�/��N<�`ǧ]�#����s��wZ����^��jյ�pW��A���Al$֎��r����ʏR�MVUj�`۠���eU������fDl��dHExY=���� \�R�FH΃\�hF��&e�|���7*�2$�e������d~�UY�����1Rb�����hd��jGDW0�.Fm�",d�<*��Ѐ߯	c���Ԡ��h�����	�ׂ���lѾ�ft�h�뾹ӌ�ƶN,����O#���~$߹�x�����'�N��[&�-o�K�,�Z�w�ٰ�L��Y����;K'��Bq��:|�����u��"82�|Ra�PK�|f�;2���Zzi�>��R��,�%cf��.���.k�c�T�K��N�U����/H�E��6�>o��I���h���Ǿs���r��b�_B�8���T���k9������#�}͵1����{0��Q�ܺ����Q�N�l�;d��ܵG�����a�p���=$(��Q/a=��XEI6m��{ߦs�G�i���U��.����)�fB__���l�M�q��ψ"����M�4���6���H�����,$��O[�̳�t~�?��,�튒`���@�0�ZN��5��/%j�}���S��Lo-�'3�h�кD���W9м���^nL�W�W=��mѡ�Y��t�M�K���(F��Eq��Ta����X�=��Y9h/y�;as�@8����޼=X@Z�����k�t��91e��5���D<Y�NFd�=հ%5ȳ��<�ΒѿÊ��/�5���$Z�o�@_8�0L�s��}>���v0��z�❦X�1��;��7��\�$�-�|ғ_��Q�5 ���+�d}hG�"�ER&�	�E\��em�O�;���c�����3կ'>z܏��4�`� �TY6~^��� mR��I�ˏx�UI����)E�̊�,~��k�1�qB/��2���r��!%��nV����31y]�s�kt���([���^���k�����	�I�ɜ�̝/���|I���g��X��Y7��&�+�5�$fA`�$kD�x.��ɝ���z7}�s�a�@���O��/z��@9�tl�Az�.L���I5(z�`�_T��n�t Ǯ�҆Z�1D�{�̈́;o}@��IG�fvT�}�-ߖ�4uǆ!|�P3��Q��n������'Ʀ�����iqQ�-<)��F:�Vnc�G��b���'��,ğRC;�vϢ|�-����7��:j�~� ����Uˈ�^���GlT�0���K5DY��N|P�r]kҟ?�����%���������<f��h�[Ŋ͸�/b&�"|uU�؞�ś0S���gr��Ƌ�24BR�����y�_'��$w��)t����JL�j-r	T���fV +�U��Y}����)?,!.���"<0����ӧ�L���9�3��Ud�4�����t�#�H�2m�����ý��q��9��\B�Vv���U�[�;K��J�V��u9yFSN@9Ю(�fe�����cL>��P;�US���
g�����x�Hj>�׌cSVS|'
�s�F��f��SX~��=tnY�E��������qD�rC���ϗ��}Ȏt���%^s�ʕ���A�.u�<����ۻ�!'���A{�d
���v��:��� �CF�crԍO^K7׽��|�$Շ�yq���ؒ| �na��IϞ��Z���9��F��J#e*_�_�Z�?��%u����T�j9�c��3,������9���_�y�W
����G�Q�&�ƙ<��w��ʓj�1*u��'d{���dc����8�s'T�F8ku���׉/�cV-{���V(3MbBjP���������gt�3F��+#։u���ՄVV��D�bW��;l6�L��`�"rg���usJB�2��:��5�hC�(�~;�C/[��X��� $���0�.�JjkF���E�e/���1�3q�1lQ�i�^�G_�%�Z�X��bwƎ�����2(;/�'r	�$�@Et��ZӉ��v�A&� ̵Yn,[��\�B���~��v3^ޣ0�����{�P��:-R��VGВMîd>\Pv�C���0{��޳�fΪJ5T�K�Ayb�<s�w3��T���1&�_�7����-s�O��5��K��NP]����̸>�֟�I4� �����3p�k���8���#�#��5f�3H}a/$�$ġ����&��d��{8�z�����������Ǔ
��S�tj�6(������������Iۓ�9�
��m���y���I�q�}w�<6����\B���c)2l��>`�p������>��<�cܐ��-��F!) EB�������W@u�'��EQ^��	ګ���3�����,҇��z���R!����?��MZ��)�4/Ӓ�x��A���L�P��۩����k���C
ddئ��>#*��$�9�wP�.*��6*@�-'��F&F�%���lAgB�ξ E�͉VɎ�'ۻ��,C�ko�E�9�r?A�e�z�I���G��#p���/צ���Wp�A��-Q����YĦ��"��8���H�[�-����4��ȡ<��G�Fm�F]}c����G,8����g�@�f��l2��V�u/\meQ=��Ni��Y��i�a-�H����(���Y;��ia?�]�ac:�.��㯵��"����)�u�	0R� �E�/'h�;��iX^�r��LY���snǰe:�7��?y�X�/���.큖YSs�}�Kc�
Bw����<Db�2�S!-C1��r�ڙO�hU�J�`n`��5&.�gb���0����yz2(�� 5�uL<@��9�,Jm�--��^�/izw-h��Et���23"���/�Ĩ���d����b%z��V���5��O��y`���\�Gi�I@G���=.���L<O�߭A�Q��,�樚���<^Ҽ��#�!{|����]3�-� �(M��:��;B���0�C(�h���'�$Op̽�&�e�D��Md�������kr��+��M������l�^��kr���c�܃[)��N�0�^R8"�-@�s[b>�H��u	M�bLj��n{K�Ya;WѬ���@q�9�֐��a��{�@0��[��m��i��)q�r��u�	j�~4�iۨ2�|���:O�Ű��=׊{�Tҝ����^�
�񞶇[��q��n�})34�qz��N�UI�}	�ˤX���U�D~�oM`LG�< G��K��x��-�F˷"V൶��UH9 ���0�hNx�z�cV�9�"����t[1Е��N5M�+W� kM�����)�,?ƿČ�v�W�6���:�ܶ����3?�Y��!��9�?�+��zg[�x�@u��,��H��r���vƩ�釶��O×Zf6%4ۃVM�R��X\sVg�Fu��z_�	O��.����;���:3�:*(�U�'�f,�0EH��3��M�y��L�N��]��M����A)�T��̳��**���T��pG�6ygO�:���g��NF�H�����6�#߶�nz��)V��ov*��+~$F~�
>/�]f9m=3⸈[5�QS�:%p�����b^/���j�g����]wP�D�D�2�4ω���h�O��KZl5�U����LzI�CA��~4�e.��S �\�N�V�H��ɬ�� ���a9�M����5�!�}�S����w�`�c��5��dn�lW�P)����:/�R�R(���g���g	7�F굿`�����x ���/F^��~Q~�qk�т���O�s�=�7m���֭9�����i��A���N���|E���S�_�Ɋ!�<ȧ�7����f��$�<7l���x��Ij�ʽ��C.�|_��_CV���0�N���9|���_��c��]�AA��%F_����Bt��@����@4j��ɑO�#��k%x���!�Wd��r�0EW�̞��v4���b�1���b�ymGĿK�x��2J�XL?������/B����r�}���Jby�4u'c�5ө�(K���� 􆕄����-۔ξ��M���k��JQ����{��nl/<q�����50�0�7�'A�3��0�6Rk@9��O��u��(gC���'�I��Q�4���Yj��H<q���*Pؘe��W�MrZ}�ʥ����W�����N���A������{R�(sB*�r�7Z=.j�����j���o^�q���&KIV��ׯ�����4(�E�-�V��sßH�k*�6ʉ��HJJ��
�Um���,4�E%�pk�NI�.�+�����O�8[��7��b"�lFLG`ln�/�=NE��n��d_?�}�1������H��P
iS�,��̄�@�1���*f�Ӟ���|���Cy�w���#<���lV�>��d ?��B%lHg����nх��#�g]���h���p:9�I���sk��5��A�\�VD��6�i�S�݀�L���@9���7i�,�K���p�p��A���H���x�W?6^��{�����H��H4q���ks�ĤdFD��ͨEu)�^ӷdׇ��@<����f�v�B����R�M�v~�R͸�|��Bb�����8��k�EaPA�� 3M��[��H}���� C��z6X�d���n�?!et4��\s}�5��ʭ�ŷJU��F~������mØ�2hO��,�D߈�ԬO6f���?Q@hJ�\ߡ4�p���^���Kz�t0��T������������әJ��W�m�h@q]�x�?���K=�z��#&�H�M�\
�C����a�J���b���d���@�vQ��!�9�9��EjUC&Q���䌅n�A=��,�e��J�׆�3?)q��`��������)83T��=���H�;?h�,m#+����w�W��*n` u��숊1��ZT��<p&FLe�F��W8�ɣ��	��1<*����V3�6�^�R�Z�I�gYn��eNq��H���91j����ϊ�"'ab{���Ħi%18�i�^pjߊüO�N�����u�-Ԋ�s;�غ��z��A����V�蝽Q>&;���&�=�R�� ��l-�YQ�Z�� �S�� H�:�O-�\o�ro��O�8�
�V �Q4�Y̌~��w�B��+~�Ds%����R���x}�D�tr}���#���,���a������M�x<!	��10�6���/�ؒ�?F�凉ܿ鎋Sn.+�y�����Z3Gw�v���$��8����fL�l���P$�o�i��m�U\6 ��44��0���>�4���JM��|�)Ɯ�{���)z�o�Q徸g��(�y ����Oq�y��G g#`�i��f�}�'�l�9Ġc�I�@�;�#�
�X�T��9��h�����Ҁ!�����g�ya)�[S�`�cF�5W�w�5Ӎ�n<�Oo�ĂwMݕ:`F��5��>	s6�wE�5�{��Ck{]S��:��~]!p	���z/ ���p(�:U$@���۫72w�?�����iͪ�7����;P�E��|�k9�$�+�2���}�Q��o��ƪ�[����,�Ix����6����	KZ��(�8?îz$@��dS`%9��I�sz�d��K���Q�G�ƑT��g�K�i=|
Y�{tZ���b���a['څP��h�z�L����m�蓒)��Fj��kdh�7���3���B�3w��������?����@�)*Z�WtNb��ٛ�Zw��;ʹ�o�l��p�u65��8|c>qۘ"�<	�����i���krw����qAPÈe���?��z�,N�}4D���˘�b�:���]�Ozl�hɢ��K<�,��S�=�]��Re��&������!1�.t���V���T�[%�h��$�VH��X�&B`����7�vD���J,5��>�1��A��3�F9� ��Քj�#G�=ro�f�C��lp��JY/�ԸqҲ�4����{�v����6zْ�t��h�=tK����V��׭P��w@�BҵϰC`�s��ş�9K[�nB�G��G���M���:���O�Tp��R �;�U3�����A�<�	���̫�J�R����qof�ϑ��@�G�=�	H�k����W`{��Q1���f�}�.��\p�C:���,��0k)�5@�_n���O��%�y���ς�f�
s��N�k^s�v�b�IaoS��x��_���R��Q��R���wx���CB��T`6�!�n�w`H�ܚ�M9�]��.gXn�����B�*�z���I��'��_`�M۸��&P�m��{�f�O��0����#�ל8�� 2���-k�G8��y5�<�_�=��/�
B�Y�b��c�\e���"�)j6�x+��ʅ�
��z���8<:����XM"�����0gE���a�����2�<��H�i��^	 �;e��<g�yȺ���U댳��>���q�-6p}_�ۨ��g`IA�Hv��GK�_�s��h,A�f8b��8D�ٚi�EBA�iU����p���e����v:��ӳeT�#��b�sn�6�-��P�y�ܯ��ix��k�x����Y�#P�n�Ρyő�єgb��r+��6�$�5?,����i`�^��<��[�`
H��JY�Y�.S���:4�F�W���ʈm���*I��q߬�%W��Y�ĸ����Q�h�0��>��ѫ^f��5�����nw"���$ �L�����s��j
>���+��"�b&��,i؇=ĹKVC#��0\s��(�T��R�>�&@�t����b~@#�v)�����_�5��.|��¦��&�xy���Wu��N�e��fh�}�St۴�bϡq�5�|"a��Ig*���}ΌSJ֭G��A��1v\`�����O�4��[�/���]`�ΙB��|$����C� �-�����ҡ^��Uoh[����bڞ�:���_������f��m$��24��enH�(I����F����j��"
\c2����gPt|�fj��׶�떐��!h�:�,�I-�/��jq�H(�N�6�ZsxM�[�?�mж�9�h��m�����.)����� ���4��?O�~У�-�����P�y8h�"c�̓��<��xț�{Q����������rP�nO~u.�f�5lӛ�k���eCR��-T���/. �i�|, j'�Q:�J������X���.�4��Z�����F��>�	uw���}��x�+��ʒ2B��0�R�.d{�Pbc|������*e���r���/���2L�e��`S�ʷ� +���jxa!�ajCK�.�A�B�S�r��'P��
����9�yx�E�
���jlm�m��Uf������dzg?�I����y�yMבP�t���1���j��g4��oF��7閪��W�&���n g�s�:ۅ�3�f�z�@D�kX�}�g�P�w�Ao!V��A��#�]o)�<�Ֆ�'d��m�_A̔E�U$�<�r�U(J�"u���s{�G�d+�A)p'��A��>�ĭ��;����X�d���4G�[�I�����/?��z���F�>���K����FR��~[����q�c��A=��.�S갼y1Ez��R��o?{����N ��٦�����L��Oky�#�9��1ǭ�،'1��u�7W�,6��5	�k���YXϑtR�L��%E:�5괙z��M�޻ )��J���SD�c���y�U��}�� f�Jg�وu��N�]���c	&uE�l��-�9��iʟ��y�v糾��@Y�Q�|�*ڛ��U3���
_,��r^܇z¹��)l-E5FO��Iم ����ɸ��d+����4��_���D/�G�.!�M�1�!�t B��h�s��#
�jn+�C��B�-���5S�Bڈ�Oxl�s��󰘅}�d�b�Z'}�?�AG#|��>g'e<����!��e<�v���Nѣݡ�f(��!��e�%�LH�Fl����^�-@�T2�V�T횞�ޠ��S������3�/��˦e�CMF���.Tړ<4CLq��|^Sri�\��8�AKh}�kFB���.�BԮC��]"��q����C�����T�$����ߵ[��F����|�-�x��أDmD8/�~�\l;*����6;_��1����ɨ����z�vi��H}���%����x����.�3ՖN\۫Z|1������No��x��\fN>��~�l��M(F��s���;��n�.=���󸘦�q<��IcH���nl��z���n�(���`�RM�s��M����ߜ�hb£��SB�9�jM��А�'�oCO��"H�ѵ$�뀞�~�;O�G:~��� ��H;�z]��t�Q�L�n�>����1
2�p��Nn��X+s{���Vn���� ��j�,i�g����b:w���89$/8a�>�W���[��I�6���߻Z����i�u<���gS*`^(-��]�}��l�S�~��Ѧ�GN�˨[{ѕ)��,L�� ��),%^x$G�unbK� A���;��*�mb��\�`L$	�j�LS-� �p���>:�؞v���i�L�(��Z���e�@�/FI��M-�Mp^�c�^�;����qa�a�K&�����-�>d����6���� ?XZ?\2�w9
���� �� ό[�Iܞ[��+�O?o�z�V�d ��1�KZɵ�j�����"��|�Vw���k�cl��w�]�����V\���>���)=B�Ūd&\ o����0Y�J��+?hzKSq/2uᳱQ�|l;bF
PS�ֲ~�b�'�C���kL�ǻs�/޽k_�~�ŗJq�����;���N��0J��e�Zx�їx��#C��H�����Q_�a�1&�f1d����$����a�i��G�|�}�C���=|��+�/�-�Lہ�lUК	�$T�Q��fܨ�RYy�ZR�޲Ya����g=BБ����x�}�Q+"�W,S��c%~k�_;b-���t*�A����-4�R.5��
�Q���L��8�dG�J���Њ~@��z~��1̥JdxE� ?- �P1 >���`&�q/���B�c~�����C��3̯���Gk���s��)`�+g�-y�t��7�M�]�?A�]t.��s�IQ6�pb�4�ܭ��90�=бZ��OА��)aq) /�����t��m��~��x�`�LŽpXMh�MD7�K�ؼ#V!+��\�sBz�c>�Z��#�a�"&��`�E�՝���"M� ���Zڋ���V������1'�ɞ�t�+��Ɩ~s�2+��Z�%�+�yH�U��?��ھ�n��(#/J��hk7�{~pԼ Τ��O���ݬ�-e����UoU���*�Yŏ�őN[�F/q��y���X�6�Y.�1��Sqz��*�3���a(~����^s�儼<>����%�%�K�6 �$�����Y�[�ԻEMݧ��E��� Nv��z"�X���d�
��x�I��A�@�b����,�o���
��!�G��b
��ai �u[��D�{p��������s�� 
w�J
��y:U�P�_�dj6f�F�a���H(Rz��_��XA�{,�3ʑ��E��,k��w��)�G(��[7=�ڌ:���%W�r��`�ӈle}�*�H�1
x���b�?>�JX��m#h;��ێ�;0O.�7B ��q�=#⿫��H�^�$����G�3̈.��VL3�l�ι����}9V�T΂Z�-M^un@r�G�u�v�N�E#�߀kH$��U�D8����2B�P������ 7�`}�tU��[eE}�<h�U��^X*5R-�y��]�BuNS�O����*F��[�>xT�*��J���_4S~�	��MV�v�e�c�|E�&����_�z�����J�i��"�d� ��'����'��H�j�9~�v����_��DU�B��:�,��0v6��Y������	�n�;ċL���2KT:
��j-��A;�<Py*xR��m]���#�c �q���vu�3s�aUb��*�ݢ�;Yc���R���{��[���5�ΞP���~�2B�+�%�̯����B脑��g�}���#*ʀ��G穫�a�����Zd����Jp�@0����\m��C��C}C���Q��챈$��tk���G$R� ���N��%�'�'�b�g�tSB�1g�����Q�l�e�8���5��$}����}�p0G��eܤg-}�F�Пė���f��׫��¿��+X7�{�)�$^g�T�����X����ؓz����4A�F<O�)�z��N��w�5�b(�0pUk}��&��;*���7�s�[����ēJ���A)9a�Ҳ�A��~�����58(���d���9id�m�	�˄�V�ڳ��3o�:�J����j�IC^V�m,��clS��k���4/u���R�G`��������Jk�v������a��+B�	��"o1��w�q8 ����VԨL.gm�����nhj�@N�v_�<_��:G�I�F��pi9��;i�s�s�-���J��#`�ND>���9���vM�Р����k5��=g����tt�:9���1��;����[Ϣ��К�����-8�wQ���cSQ����(�3K۳��B1�=_���b����j,�3U�I���Ck�i�Pe#��7�9,��5��6�_ ��5�͖o� <��B�k��TI�=d	�p��Iv���P��ol�nP&ӿ���Y�3�2_�$�PnYqL`
��h�A.���ю8�`���C^0�GQ�[���K�r��7���aH�J
#c��I�p�����
������c@���5���[� dP�F=6��ў�P�lJv�aǽ��u�_�����w����pJ�+�$-je�v����e�(Q�Q�d~���&������!{�ލ9�RWUB�%�������5��$[ y{����?��?m�e*��� F��
W��}V��d�@o�uN`�T1V��PB��D!�	"�����!��g2UAR��e!Dj7����]Rݖ�j~�P�	'u��_ĩq���Ut�u��a�_c,$�L��Ʌ�pѯ�ݚ)�v�e*w�iC#!Ԟ:�YƑj���C��9-���b�r�@��5�T�s��i�T$� �q� g ,}��3H�x�j���M��;�n�Ҹ�TZ��<g��s��a�Y-����]�AIyj�+�u#��Ml��d#D�c�4�
A�f;5uw`ܮ�"�+�G[8p���>2��o�{0��X��p1a �_5m����	���K�A8�{p�EP�=:��S����~ t,����m�'K��(�h>J���$z�7�CQZd�O��C&q�5,;9a��!�8X�K�~vg����1zdW�%#�����/�=+1�BHQ�8����ɣ���iY��`^�o@����ⲿ�n����9�������$=J�U�H�B�KjG�m��-Z����I��s����>�@�/S�[!)@輺A^��]�A�rFK��!k�]�NǾ$a����d��<�y��:�-��w���bO��M�O׺�t{��GIc:~%`e��`{n�4���kt4��ؾ��[���ɻ������;0�N���PUD6֧�����9���`.m��fn�נ�b%�S����B�*@���k��l�r�&��?�X��LUr0(�r���nia�ސw�N�Pzq_R��Q:i�N�]H��	wr���e]3�h~�V���	`�Rv��<�&�F���<1�u���uR Er���[�6��X#�+*s��!�ҞᚄE�����v�_BAp<�o	��LL�Q�A�����'����i��u{a�Ud��� ��O�4\Y_�3e��2�1��¤qAw���?c��"���fct�@Q��;oVnU�:�>�6��DM�Lfv�|oܰ`�>
d���3���;-�g��ب`�j��A!|���뤽jN����L��dã�p>->!�������b/h�0��/�yU�]���F42r8���$���C��U���%��:�A��8�'�����������emr����R�H+�8�"\p?A2c�,�r�Z\���S����W_<>���,ya�vÅI����ӑ�3�T�Mgeʔ�7d��QG5�L.��1c-�Z�"vQBJ�{�r6o޺��Z�'�	�˾����]dG;F���� �~76G��ޓr+�J,G�!?����k��x���� s�9'gz*u���v睎��C�\I���Ȅ��v�~�����~�6�d ���NΚڄ�m�`G%A�«�� �
�םl�w����@F=^�U���"]��|�N�����/Hh�CF��9�"ӕ���Ӳ����g�vd��.��Z �dat�Bl���H,��	��(@��t\pn�� �e>ɬ+l}a=�kt�� �	r*�~TeV���y��3�R����7\-�S����چ�����r%P��:�����Za�)I�bHo��K-��G�~$�c�rW���m���HԺ��Le�����ߋ��CeTԟ�!��T���^X�����__�>
5}��z���-W��8��C��X�29n���t���h܌<�f1��D^}�	L��(?��Z�����V�`y�Q)nz��y�	��ż
���x��Ԏ���:]AK����4q������(��X�)$���Ώa����ۖLvzQl��ֹw��K�/�P�XD?�u@*\��d�V�%p&���	T�DPՠ�6��^T`��C�c��ۙ:Q�2����Q#�(n�ɷ{����Q]Ԡ�=�)J � �Pl �|2aé�e5*�&�����$��)F�C>S�m��d ?����l�C�<*��\�}��w��*�I�,AǾ�.������)�q�VXi��$��aQ��T��#�GF"򲣥pC���Ow�j�\.5��7��2¾6�����q����� {��R큡2|�f�(�A��(M1�U:��0(`��#���m��b&���ѥI;���-dԣ���ά4�B⻶AႻـ 3���У6cM�G��*�>��4��G�?�"��(���+���
e�m�Wk�� ��S��/c1�\���"�<��l,+�H�UÂ{�F���7����7��������)>Z�l�Z,1	�2�ʃY.ڧ�'�ͳG�%��نw[�iH�&8��ja:��.�����6��JX�Ix@ß
�֠_1RjFp��oH:�!�a��)�xQ4B�k�ɍE̸�B��΂���c�[:����4��s�c�~�)���[d�_΂����6n섘{#�/%<���5�t����l��B�S0�s9��CFy���@��U��I}j4��&@7#'M<�����)F�!����Y�ϮO�|��KW<������W�O�f$�����!�FA��Usz�Ê�����EZq��'3"��0�M��=ѽ��*-*�oe��)S�ψ�&��2������U�q�V�4��� X9� PD��,j���>e��%�HG�k�N��Fr�W9���Zi����ˏ����X��O�c�b8�����v�W�f0*Z��>��~j/ 
BM=U�|D�'�g��)Ί@������"��e鯆?���
�|e�u]l-H�)�s=����X�����wD��L�����FcD�� ������֋���\,0w�^��O�?�dl�Y�r%�4������ ��V�A(%�!1[�1�8N�t��T�� \�P��+�zNz�Br��c��4#`P�Dݗ���k�Ա��Z�J�!��y���͓���dB��:-,��'$�m�O�&��0���9�(i
��
��G���=0G>e��J4�?��/��P���jñ%/���W���Pa�@pk�!��,��ah�n(�~" �Qdr�g�צ �9�s���&��_ԍ�M^,J�������$9D!y�[��������d�pz@h�`�5�`Y��T-Aa���xky�Ƣux�2nOD�����ߖc��
���f���`_�M. ��v��yY���8���@�{��|��(�zV��z��͒B�~���DQ�����R�wپ�4T}����b���瞤�~��&1���aӸ����KM�zA0�
Lś�y�Ṁ�Fē��-,\�mxyt(ߏ/�H�}���C�n�V챙��r�
%Dܟ��X��-�L\K����s;rA����q=D����e>��rF�i��ײ5��D�F�ؿ/e؋[������c����U�k��rW�0|H�����"�@�f�n�bD,c�׏.��/�W+��i��/�F+�gB�Ns}��)�=L��ԅT���Egy��2�i�O�"?�8��q���O*��!�-�H��i��
Ǉh���K�13Q���f*�} :Q^~'��G��^Ӵ5j��>�? z����4&a�����T�8[M'Iv`����`S7h����e���%��͈�[U�2�ⓡ X�Jp�+�4�X%%�,ّ}do�7�%&\���=Ӽ���JB�M� ��܉J�U�[�q��j������ ��^tM��/�%&��n�i�~���I������H�ڷO<d���"�A0p<�*'6���
-����V��,_�>i��p>�Zud��蚅
K���M<�x����w�*�aZ!t �S�~�����~�F�.������t�@U��%�G�V����0�=ۉ��h�7�����=,Z3�&	H�k�!�>^���m1�6) �aO�|�N���S���_V�C�Pg�������^��`���Ս�����BD�EoPY�j�SG�1�p<�UV�`r1像��t�쥇��܈�2����C�/��Pj�P� ��o%��?ڝ&�$��I*!�e����vI$�Hxk	8ܷ����S8ZH�
��4k>�HRQ��Ru=s-�v�N��Ӂ��1U���.T!���q_RU��הBG/d�W:�e��-�Ŏ��͏$��r�5�ތ�(���9v`�a0*��{���k� �6n13���z�,;@��
?��¤FP%��ggݓU�\��rzsϲׇS/��w2݂��t��\����X��B�0�=Q�i�`��ͧ#W�3x�PY�,��(�@5*d���c�\t�&�p]ȋ�p��b���>g��7A->�nx�(nR���{�<���$�b�kh#,js��Ƕ��6�^���H#�$���/�XU)Ģ\��/�3��?���u���?���]�ӴX�4��qWL4�s3��&�9�N4PG�}�{4�j���cxH�ჰ�_\�r��7(�]4��p�=�eX�w`Y���:��X�(�7'�g n�M-��j���!�ҏ4��Ţ��sJ$���U�G�%=Oa���{�X��i�xЂu��q���i������\ǈ�f���M���үf�x]Ь��kO}YKAm����~�W�XHƝ��,=4�'w�R@:��aH��V6�	Y҈�ƬD1�|>����X5���m�֦�B�c'!����pɣ�Vi"!S�ܩ�� ����r��@L�t.��^��s�zD��V~����yaC���W�+'�1�Q0�(C�)|U��&~n��j�nH5�qN���?��/����L>Z�<!�Ɠ9A��e5�i=#�m稉pe�\rt�0�K<=�:Ќ:�d;����ݶ�H	�Z2���LSZ��p��d�Ż�d�T5�s}?����0
."<~zw���B��_"M,�
�L�&·����5����>��=:B�X�_C��i7�O�.,7�����i$L���@���~9�S��5�ZNM��ODOv�3�h�������-!氆̞_5"�#� �G� d��IPȆ9�<�|����m�V������z!��z���;�2�F~�Ӣ���^OU5sv)�����-�RW���3a���zr�x��3�j<���J��Rum���~D�*+f�6�?gP0��P�A�
_:����5;"�4 �2J<�p����F`�qfX�a��3�	�!��2*�)��5��2r`J�##��ɺ�:�p Z3�������	7zWY���B���˽n6�s@ר���o����G?�H/k��ѡZA�;��/$1&��ʶG�����p!0Vv�d��Y0�A*c7�n��6(�(���|���ﰳ�DZ�	��/�C��ڡ4����������祰�+>�64i�) ��wGV�՘7�{m�f�=�����
� ��K
��QeLǍ��V��kIr���dI��BC��մ�R�����������3�����MlQD7:- �~c��5����2�\3��=m��Nj��J{�ns_M}�#2tf7��W#TE�=gSGpU�L�X
J`.,GP��� ��ٿ�z�/�� z��G�Z�0���T�Ax}��b�J����?:Q3�nX�Ec�гw�5�_�Wl�nU��'��,��S#m�d�6C^Tx���mE�N���z��#�}�̭e��Wt�V����Y�(61�=��apld�^����q��K�+5GF~{�yV����(`������N���|�lA�/��riÈq���p��l
���&�hT���K-=N��=|����h$)��)�~�[�;{U\�{c�J#�^�Zs�"�(Gi�R�w��>�[6Э�H8%U�E�/�n���j=�5_��7�tcwM�ï�Mh�M�ԱF�tql���`!�x�[O���WO���{f��j�OKH,ޓ�f�������Οc�fxq�`�"@�9�+��&�Fą���(���S}��g?�]���b���j�V�w�<$��/���o3R��N��,��EC*t��kۮ��be�_)kifI�4r����c�kз��$����6J;�2;&�ǔm�Cy&�r"�"�����
���I��M�xŏ;op����Ԋ4��=7���g�v�'�x���G�<���O��;G�#B:,�y1���WE�S?*睾�!�E�$Nb�[��Tqw����|i���귥|��2 ͧ�+����ή~ !�n���Vq�mU&fCk�%�տ ��ø���"y�t�h|j�P�&�	Z�H-$�9O�Y꡾x�fi;ûe^[`�����,>0�u�HX�G:O����s�Q�ի@�R�n�?���v�)���8l�.�-Ƥ�����=*ǉ�3/zO]@nCe8t��ވ$�#�)�w��hտ%~���?
����M	9s1�Q�&��͸�'�	9_��1�v�O�q��Q.[T���<z�۾�[@�J�SzL
@u[��
[����5��IGj��`<���� $ 0��f���q��2�I^���g��ރ�f#o�5?<R���t�$�^���̬�4�]fx��Z��&BO���X-�#���~��f)۲��5e_6�9/�O��h��2/�6�����k��-h^�%��?Luv�����D��P�KCur�����g���A���+���'��I�9���p2�����}�O�fm}�?ꩋ��3ژ���1E3z���x��U|y��ɂ�""Φ�\�p���|qQ��[��!0ݺ��	��z�c4pz�v����B��[^�d��Zx8��
o5�#��	u����"���[ْi��q�Rqk�|�m�"��­ab R������0n��3O3��0	���;��������ژ@5&�g�_m��&�2�[��;+�@Z�h�6*�g(����������;F&��}�&����E\�f\6�1�
h��¡�yQ�qF��체����Ý�9!�튂����'j^�lt,0�y�z�U�2y�1O+�.38�$,�P��g�M5�˹�'H���%����qJ�����O�4U��Uҟ���<������L����Z��Q�T�g(6i�院r���+����C��� ����L������Q��Xm*�(嗨Ǭ�{�!lO[
��#f�.C��~�,c�[�'LdS��Y��%Y�D�f��."��?#pv���Z�+@���6����8�pY;3��`�=��J�yj��^��㱌�!K, 4��j��<�}=唂)���Q����G�Py]�tS��J4�*Q��Q|B�K��F*Z�3+Z��9���i�9�#){8Hdy߱ε�ڌ��h�D���[���|���
�-�*sb~e�S��@?�Pz�Q�J[8����t�R�o�r���r|7��
ʉa=�Xp��64���{�|�}T�~����I^���{>��9��"���<�u]����
��f�ތ�4���0�G�a�j�H�U���&'�٬ףԜwT�#c߮:�8[J��m�·�˝w�Ȑg�*N��l�s��;����c;?戌ӷնI��m��B��!�?f���ގ9�	�_R�`ʯ�O73���	T%.�����,��&�x~�C?�	�(���:mFB�]D�S�^%%���o����(���PV���k�G�@'��_#_v�~XR"IX�����vO��I.�d��u���!z�'���������sK08braZ/����3���10�V?����$&�2�1�̃˖/.�o�W�
eM��L+��0-���Ie�����qC�'THrd�)XjG���A�M��^sW����:��Q�rQ;DߌxQ�''�8Pb�ؐ�>9U9���L���y�^A.TD���~�N��.�#e/`ڙ=Z�S�
��l��ؤhZ_2���e�i���b"qR?K�j���fr`c��*h���C�R�oG�O����4���AJ��kS��h)��Z幰E�Ş���9Y��"9ua֬f�=��BD��Ǥ�O���<�e�O��i5���6��y��9?��S�� w���Ͼ�W� 6��%I��1--^����ɳ�w^j�h�����N��ԣGmU=qPv��N䃳 ��:�:�q��N� 7W��S�S�1l��uSW;��`��J�8�a�!r��"B�9�]�m#�J��c��-���k)#��s>_;�Q\=�T)P<���Q�1�V���g.7�Z��"��N���q\�B���C�UTcW�o'�Gd���h{bV�	��M�����m�ԇ�9�_nAE�5Oށ�4�X���C"J̅����* �3�������|�#���B������� �W�ԴvU�-Q��0�Oyϯ�v�6�����k*����4��(	mfڷ�n�Ձ�Ң�6w�S��@����$��ޗِ���	?���/��7����lPz&:���3�l��O�U6(�>�g'�V������X-������S�^(	_��)�[C�]P�
��D�hY�y���Aؕr�HUv�E�����?�9���4#���L ����Y�&k�M]�@�� ���$�s� Ą�E���y\�a_�1�y�$(�-5"������O��gYS\X|b���`�m�?���)��t�@y����ͮ-7��v5��c�a�]��H ��O�K�Pgn�H�og.�0hFPG�ۺ=��w-6䛶�p�����FsGJ��hMK%%)� [��aG<�
ٵB�`�����Nx
t$i���ڽEn�-י�]87ֹ���?&�;�.�?�a�D��q�:�u�9�N8��O܇�}-����ܘ�՘<���Z}?z�H� %;��r�����2�ƫUd�P�X��$��;��� f������?L�׈�]Hy7�-סqI
r�z����U����SE���� f�-��K]ㅮ�1%"Ir����)B먟�~&-�Y]lp�S�i�wZ�t�ᓵ���*�<M2����e�át�}��>'�a�gs�A��2�6�t����FhL��x`]F�\���H��H�V�j��?Z8�I0Qжl%f2���t)�Y��ʹUq`�tKj����!�r���kh�D`� `B��U{���/U4�:B7,GF\�	LWT-���.!T�u��v5��M�/ZX-CU����R��yU2�ث�P��{	���Ɓ�0y�w�6$lԿ�`��*%�R���}����� �59f�K-��� K�ÑzpI��֥�*<˭�w׉���烩�tП��b�P�,n�=Ul�վk*i���H���:��v!�/��e��zrjG����`��"x��Q���ek�����Ț�����^�������q�	~3!tW�m���Cܢ�k��1���ߦ'):,�'�����S��X������K��9�=<��e#& txt�J��q�F�W�(�j���и���f�"8�Z�G�ʭ�ɻ����5>���=�42k�z�!�i��M�g�*_%����<V�2.u���n��&����r�|Hı��`���Z�c(W��5U<��-�;�	 J~*����d��kv�}�)f�+"(ob�I�K�D�k
����^����s�8��_��da��q�R<r#a�;�^R��BQ`z�nQ�b:�]C�l���u�	�5nCͽ��\�Wr|��I}��jS�Vg���w���LC�����W�j��x�x�\�$�4vzG�h�A�AzA5�(с�^暸�(�
��c���R��L����m���MR�`]��ƫp�_&���Z�Mx2E�KH�^�[�X҃N׵�8_\[�ݞT��B�.�8ґTե�� ��YS���_���D`��C_ciS�%!�"��e�Rv�ILʡ���&d�v��x��"�\N)�>�2�1��J��Ap��>�D�Ȳg�o�ن��ᓽKyR��i�'�Kκe+,��X��ʞ���/���s��%ii�Y��H�UDH�|���0ϵ���0HrmʢU�t��:�WÐ�Ӑ�4�=nЯݎ9�DP6[9�#�^2d*��S1��85�=���(�;��\�>v��l��Iʛ���&�$�@0��A��7U�#<Nu��[��2��1��j�d��$K�:�����\^�ْ�);�$Z�Lw��������#F�%�vf��L�E�i��Ysi�=L��y������މd�8vN������;F�f�w6�-�5���ho��QJdT�C��'6h<:k�/��(�&���'� ��4Ug?QA�Bۍ����P�:uEۃH�b��
��Ѭ��j�'iv�?;��"�d;$�xp�6�K�R�M���_o�{�=�D�hn�O�|���@��K�i2�5�c��8.�E��8�iQ�H�8xy ��v�t<$hC$1gSKy��šu��~�d��Uz��gnBpSUɉ����P��|��%�c���tPy�����\,nA�`�_$�7�X÷D���(��$}�.�3�����R��"�
9���@#��C\DS�"r�X2��,��)���=����ɘZ^����*����ǳ�O�P`���M�#wk��h'�{�!���ۯ�a��}Q=����?Fv���E���t��R���E��)HЂ
p����V(`	��_E	�E�˗���A{�b�ɱ?�\͋�I�F��3��D
�ʇ�E���y\�.$a)��L��B��bPZ���)�8��oPH��4�b��c ���̽O���f�XZ�f֎;{#�R��]H�졄�fޖ�������ٷU"��I[@�Y�m�����]<�w]�Sݷ���m�-uiY�����T����Y{Y.{ELtIk��ڼ)�cn����mH,%� �I��mnAl��qe��X�a<��rsݝ1q^�Հs��K]�2�7Y��Tw�0D�3���<Ѥl-�I��̚�珗�N7`�ì�D� �Q�m�AZbWn1-�(�o�����ǐ���[Ug�x�:RB��aY�H}����L��&lS�9u�Q��i��+V+"�RJ ��0�639sÀ��(�QtC�s�A����(2�M�C��qfs��/�@�}^	Xo�ޢ�3Q��3[�d�������i/`��.�Ojd
c���E+dH1��� y��8�&�V[������RK������p3�00/�P�TŷC&����;}�;c�6�$l��yeJ���[��t�M��z}�Om=<�.����'h�;|�LP���s�]�7}K���aWä�XN[��+w���ם�&��_vL�k�KRŅC��k��6�#r9��L�!1��w��� ��vڧ��|jͭMW-?)�����ہ�k�8�B�+e ��zjld�kFT��,�s�0��G����W'"֌4�e�'�"����Q/�s ��Hņy�'�@t���u|ʊ	.b�f�4B�[A�s�m׵nL�����F{����<zP�-X��L��i`b7��.>r/+���6�����ň�~-Y��ᷙ<@�Q�Gf�*3����1O�]P�O�"�S�q�8~c�K[�_ Q�]�0����>�HrgL��I;��-��5x6�����-z
��9��'�x��8~&(��Ш��"�3�1�����	ۆ�$�Y�n[Q*��'��]s�-ٕ�a�	��ݐ��l�c��o���b�	Er4(>!��$��?7^�5�^�$��0�6�����ט�Zŭ��d�EO��YP=]鐣t�AR��:-y�4��6��8#B:����.V֠��D��RU�#O}S�F_��6�p�L/7�,Bbu�r��k���|�\&���)�IY؄�������-�x��e)G؇���Y��|�|�i8�E��̉F�TɅ��_��Izm�i����G��`��ա�i}���sV���
�<9w�k�%^�v��^�� �o��|����  A*�)"�a"�-h9�N�}��ec�@<����"�R5��4�;!s �94�Udʗ�Z��J�f2 �ّCk�Ҭ�>�lq�O�gp9j��x!�o�-y�&��+?Uzj�FǏ&K@:���"Ec��b��;�kȼ��>��/hZ`�Ts�u!,��(���4ѝ�[\����e"(f�=_T�8 ��ao�e��)��Q�R�^���\y�?����E�+�YF�_��^��f�x�SR���*���Y*u	���q�۽�4(�=�_�g{�o��'^�J��GJ�B�	3:Z7 �|\D�x?�ѳ��ӄ
�<��0�	�ym�����o~�Eʸh���r���O+(�ؠT]��f�n8r�0���U���?�����,R�Y��=�{v�]J�8W3�'����n���T���:����|��Z�TK�ѢWyqgy�����|�ӣ3! U��iwr��f����N�U^������a��U�xU1s`�3�c�l�!u�y �a4�;3P��Ϝ+ps�
Hf��l�;���pN���~A�s(2���r#��uǺ�'��c�?ʨ�0��e`�n� _Ʋ�q:��!�k�O�f׉�v=O~��b�;�ֺ��k?��g�/�	�z���e��e,��ْ���s<���|˕ ��80�l��\�T�hP�&�d������60C�D��y�,jӉ\7Wdx�U{�?ގ�NW4O��l��$#A�4����Mٖ,�Y������A 4�1����Ei&`��ۏ{���r�M���
�����驀��[Ij
������B���Jf9��+�k;O9}Eik&кq�\&G�]݆���O�J$���5";|��g�vX,�/�i|��
P.�k9�7p��r~�)��?E��A8�vryx�� i��\�>��̳'���R��W�{�Z���1�.VT?H�B�1u�gѵ�;'��� X���w��=�r�Z?q/��7��3ǖ�[ĭ|f\��c R�0�����ƣ�Mf �G��^��*+��ށ��z_э�#DUC�ƾ�ֶ�A;.=���~�	s?���o� Ɨ9u�su=�]�ˉ�gr0��v����:����dS;t ��q�
�,)-�q�T�]�Y_C�)�h�mLu�{����H��2��DqA�2��
�x����U��>Mp��c��2����n�.��bXNr�V삽U�ЋLL*���t��`W~��s�)�|����כ��M�_��	����g/ҧA��z׍C����r���:�#��&��(+�'f�|/a�i���:�8�7�b�+�hS�]|�k@��d��[��%�����&�Gz����S-��ڣ�WRtesa�t�R\�D�/�ؗ���A��EF������<DTTA����c�x��ζ�V�o��[}>#�RJf�a��{WkJU��޾��N��m>K}�@|��c̓@�T���ua1��>f\i��&�4��q��OT.����*���2_��Sm��V
֎�`�	ޚ�9��TE|�{P��"o6nL�( j�;%��|� ͘���`e�����V��z8%s#��[ߡZ=�`�6�7�������Cne�I���bu�qj�E�d*8��<S	�nҜ<�w�%o O�W�=��/@j���B�^{�כ��F�''|W���P�0lkx������y-�����}8ɒ�ܐ*?���������G=d�n[΅b�+��^C~�5�۫�@�x�w��u�+CrK��>3�p�k���ox�=	W��B%B��h��m�` ���!��~|��#�9��X�j)V���/R+�:������,����1M��zTf�-���"8����^���]�	�BV�K`��W��&�`c���{=]���Ƨ)�O�3Y3k���\�O�
��V����)�	A�G�[�OJ�j m�`�Ϳ';Fm��Q/�z��p���2����r��]�ˉ{{��Y跪k��=	�P˨��� 3oC�G&D]s�[B�#<sni�<"36sO����h�:�;N�|�������Z�����N�5[ME�w5W6��a�G<:���OT����Ab%Vs�9��JMT�����X:�/#�T��1a3ae�>��ZG��!���c�´c��}+ԓl�`��Ԟg%�Uȟ�N6��g�t�ǯK��(���Ќ?��]@�fm��b�x���&Ȼ�a����
X؊�I�4��=b#�6�ѽ/9����P�)� H�J�@�q2(&W�.s��] ����#X�I�j,���zC,���9��˒Q��E^k�t�!Z�c���	���N�Dٮ1k�\���洨���o$�@/4��޺�"�'��ߔm%� ֡n��
:�/M8��I��8�&N��4������'I�m����̀�7 ���h&J1�s�}�zlJ�^�o/%�5�p[���"�[^R�s�ő��
M�E�2u�i�����gJ>+j�J�c�>���g�=X�$���-���+]�n�/�XPPԓ�/��V�qC�i�\Fj�μX1s���������z�!�馎M�HcQ���L�7ԇ��9��š��fu0^|�S��f���������_6�4ɟ���⅂��Otǉ�y��K�T$Fx&����H2��I�}g�
	|a Ԫ�W��
�u�'Z�c�:	�H���&ܿ����;~T��O�.�#��X�h����J������3�NA2�����M�Ȼ����˙���0.Ņ|)%@�ڞ؁����ʕ���,�6��V�Dѵ K?�����/���k��}[�Tȕ��R�A��b�^r��8 �RJ-Z�]��߻�i;/Qkޔ��<��l�S�X����g��?/VN��>���h��Ы6m\(P��Zk!o��{e�C���Ԝ���`���c��\�`eu���&���C��n�8v-TZ@�����Ӵ)�pjR�S�e����N{{�/�5yo�r��
�@8�2"��H��-�;˚����R��L���q��5�_+5�9��O
(zL��M�<�mr�@]Ko����j���7�y�9�s�PZP���7^�,Ŷ�ّ,�Gx�#y�$&�*���6����B:�<�׶ߦ�����0�	E �Ax����u9�MG�_��Ւ>\�^�7/��h��CI�1`qC�R��|�Ԏ�W2�li��AZsyX�ş������ |FFGȏ1'y߻�*��yOWL�F�uU/�U������b�eNa�P�HYB�J*�A�p��Fc�N+�F�)?'S��^'��5\~Y	��Ʉk�/���/��%�[�!C�hJ�2bhnm3xF��?��鼑�p�$/�Rx�7�>�<�c-f��{��d\q|J�i��¤��zv��-2�N�qZ���Y$��X��uEe�ͦs#��a[���
h2�"�����]��� j�R�M#�]��[��u�߽��mq�܅OF�8`kMܭ�e7@ 
�(�6�����C��_m,����cZ4����&�lG�һ�5bk�~�� F�=�C�щ�y*�7��T���	s�u��Y��~v\�8K���̨�H����GA�1�a}�3V�E���S�*ݰ~
�9p�z˸#��:�w�]��K) ]�n���8 �iΈ��k���7>����+t�<&��������i�Hid:ͭ��8�8%0�PK`|+B��?��)T��
��{e�%:	�*<�jkX�@z�&\J� �<_�I��<�XZ�6!�^Z�t�O�2o6N�\��J.���ڡ�p�\�Ok����)g�,4;Y��B�UU���(�M��N7�	{X�5��qճRR2����Z�<��6Ol谺���
 o(�!c0�2y,�)��C7��c����0�B�N*6� �O�o�:�=�n�A�&�f���\z _��u�/L��Mx��D�n'�D��XjL)hs�&�m���3u6`~o��ߺ���d����3n�Mgj�j<� W��=2hI�F�ATg'�*�%=:�;�+�yV����(�T	�ՙ滃$��
\����f�#�95���\rDR���b{�
�@�	Ȋr"â�Ke3�MD[gߘ��v|3>Ӓ�)�w�hG�-m�M��f�1�EaxM��F*.
�sg>T851u0��Tjv�ˆ�o"��ny�����;�f�[��|��P��l����~bZ�lAy�zf�̃��#E�$�7�MŌJŖ�N�aX b�4�\������#SH�^���e"5*���[�vw���r�r��Ǟ���4�Zv��� �{��ցkXm ���n>4Н�:����|�(��5��}`�H�M�v6m6��?�JF3������좔�߽`�~������=xR^���ݬ�ś�⹃>zH�B�&�8R
������)��L��lG�W|q0�@:�)m�M��:�L�ѝ������4�PW��]��~о$��� KlE�aYHɎ7��Ff���w")i�_���)T�z2C� :	�᧥�/>��l�x�	T��լ�2ܵ����m
Ez"�ן��F]4��AQN7��4��{yp�4��P�jw�w��J=-�Rz�W�HE��Ht�1�Q��
�9�V�y��Ǝ����Dv��M��e�=F���e�>e_:����R�+�pCgw�Y-�P>3��HO�֦ 0n@B�E�ʀ��7Jߕ��9��&
5\��3y�F��!��-2˪�����EF�F��/�����&�� ����8�Y�U)���>� &���@0۳�ȋn�b��'�L�g���d�\�����4G�X���O���rfO�(�i��� h��7�H;nc�2ҷ����]�D�p��Rq\�]���@��/������w�l���n�r5G��j�]�Pz�h넢	��%Ȏ#9]�<�(=��Y�'�;0-�kU�2�3�}"u���۹�}��#���B���������j�9�o��TT��f��5; �����W<�):� 	��[��D���k�{�wm�N�,ʥ�����F.���f���i�.���͏�sv~b��x�|}�y�-S��%yb�2,(�Lw����׹1/��ǧ^e�ǌ���8�:CjR;�:qC��˸"E��(�b���f��1Cql)�*OUP�Q831��`�k�&UJBqw��:��5<�I�}JpDֻ�7B' �X�����aY�X{�ʗYQĖ�:�/���bÂ�ۨ���������<�s� �^�c�,I�y��A<�δvrl�ΈEsZ1��fD\�K`}炂X��w�iV��YPw��5��2����1I���� ��T d����_�����K�зZ5�n[�q�tۓ�sQl�0�O�B�W3u��^���P'ռz�!�p�Ӆ�����]<}G�|���0�/���Z>�E����4|M��x�'��Ǹ��F=+�T�Yq��Z�Q80�(]�
4t�Z�5BG�*��.o���� �Տ�kK�e��ÿ�=l��4B"���;��?���R��l�����:d�3�F���ܚ�;K�ԅ�M�)ʺ�t����;���ze�_�"���جz媐2�X  )��Hɲj�d�\Qpȼ���#	iR~����&�S&���.������uKm��7Z.�ު G���m&+2����f��2�7>�;��(?�e4��t�h��.^�$yޓ���:RW�
��A���뙭�yoJ����mG�p^�ܭ����ՈAv�N߃��Ƭ��K�S����R���D�^���L���	;��Ah��{yq��`B�R�������D����uN�������
Ѵ�#E"j㡝j��DЛ���_�9
"�P���+wKm��PP���G��J�?d��HC���z�O�!��r`H�J��ϡ2�� އ�LZ���8+��ai��^�@w^KD�y"�4)�Q�p�����X�%�C���ٴ$*&u{��Yl�=j�����*9:e� �-�_�7�����*�qh�����.IÕ�R$�_��ad��q�������lU6[p;�'���t\�WJ�U�Z�=�-�Ir��C�G�r�u����?���9��Y�B�e���ߙ��x�K�.ʗ����+]�m=����hb��$	���j~�-*��_u�x������c��A/�2��,�g�o���c^`H+�AW%��A����-)�JC7�!����j[nr,V��En�UiK뤎.�oU�Y�g�������u���5�J�����#�G�+xs<*��(ϔ̐u�r��FfY6GVZ'=b
~����}���yK�VD$y ��IT�d��/,�b���?��\I�f뒄~W:�-@Q%}Sʡ�T�i><�<��&��kVǡg:�/�Y���K|�E�_���H@�(}��f{�ӈ�A`�X�r�������x�մ�
��VE�+ý��r3w�Χ@��y��q�eη��2#�%��8�xgV� �Z�:< �`��V*%���U=e���d̽�wB~���F�eLXr)��y�"�28vRP8o�릨���m<�$rz�@M溬�n�a����m���?6̨��Z�%��3�Y0��H�4��}�P�$��< ����Z�l�.����& nX���0:ٷ�p��������~�8A? ���K�r���:6����`3���˶���#������7�L4�RѴT��5���V܂nQ��	W'���9K��V�4;��:�d,�R�s#m�W8���{�L��ŹQH3g%֓�>$-v�C�U����	I��E�-Oq9g�M����i�8�Vr�<4��qEe�A���n����]������->d��ܝ�3{���3���
��#����(���\����Wz����t��*���F��D���Y}�Jͽ�h��0g"GV��<���#a�3�(dg�&0W;u�29~
մf3@beΟ�=�n� N�A5T�b�f����t�F.�_Y��q%g��X� ��~�|f�~�+�ŜLA�{<�(�͓����h���.�$P�{�mO���f&p{FGvt`0���ٖCE��Rh��JK�?��z΅�A,�+�HN[w���0�c�F"� ���Ь1%U<(/r��+Za,�H(ZĘ�ТHv+��7�zm�A�.Y�!k;"��#��!W:T���oR��t/����b($�F!���SH颾'�PԮY��&b"�M���x]�@�]j��X�����w!l7�nh]	����i%��K�$[p&�,Bg�n�k���L(�abn����%{2�'߂x�D���!�I�S�����t���5���2#��!D��jN�L�8K;�yZ2�zh�pەԚ��̓s����X�O�|'>"�0ӓ|Vaf���HnY��4,����W��<y�v�z�&�� }��rP�L>=���8̯���wQ@G�հ�� ��_=�ر��]"���i�y����s���ܝ55����J�HH��ck��<mOZ�+_`jU ��yA���CU���8�
J�Q�	O?�B��0��P���J����t�Ue�vv4G�C��v5,�`��A����rR[1<>
�*�O<���������	=�m�^D:��m��Q��G������Ԃ]�&��e��3�N�'���Ǔ�!�&r: ,�U~L<yg@��?)������r��&���ĭ6����g��X�"�*;������C�.�Ϙ4;��b�%M�ފ��{#�K��BXc�����w�%��Q�|��VL��	������.���!�9���FG�*_�J�͹�Voߖ�́�*�a$�bP4'�+AO��5�,���
��7���1�!�F�m=�s�h�]2�RH���USf�x8�e="��{,,k��M!��8�c��G�
�zi�2oD&�Š�W��ٵ�m �����lFi���t�b�%�7~�f���e����[#������JJ��	��j}��-q�ū��H��\�y��uC��|4�Ǝ�3����f���-�Xss-���
��] Q�ӄFȾ�"kL�y���H&����,�Xa��[����W�@՘.Z��J��� ��%Uf�̔�S��<vJ6��[ތF���E�&���(:��%y�t-�M�#��I�(J��A�Z>$A�E�U�d|>�kּ.񫄌@�r�r;������*t�(�pZs�VaA��������)��{�+�3�R��iS/�.�^�P#�	=)TO/�܍��)
�Lǈ�ݞ �02j�<p�NR맕�
������f�e��'�	P	�6g���Os��BW���I���M޿u�!�p��kǖO�<�$��,ŧ���	,L��,ER���"��4���:�|��%p���͚!��q���� @]R
K��M��-�?c@��M�t=$Y� ����CM�!o�4X�@Ǚ �`���`~$�F�jҀ��
��-�X"�T��2 ��J�ъ�(k��E�������s�0�8�sԤ-o"�u�{L5
���S�r�h�j����*8T
�ަԤu�r�R�`a�դ+c.5-�E_�_�MfT�q.�\Q������O'?ŏ�W�jd��#������xW�Tʠ�>�8,[�{�v�����	�t�����I~
@�(ѧ��u((�I���<�^?��&.��F0؍֢}{�@�<�>Y/\�: Jz��>���e����.�IE�#|:Awiҁ �b�Zܕ�����j�:~��̄�oI��ϻ��o�V�P��]H�����������M ��t ���`�IĨ���r�J_.roYJ55/�#��5�nrte��WJ��̨z���jb�"��;Mޘ�R��J��&����T˳LX<}��xI�Zݱ�W���+	�Q��9hD�W��D`x����jt>V2�Z�y��6�;O�T�&:�0�Ģhboй<X��r'�����׺��N�N��e�|�d%X,�����\�,QQ���H�Db[�F�z��F�l� ��A5���ʌ�Q���BR�>��a�I��lX6�)�(]T;hZ�a���xd�����W��x<n�n�Ca��;R]��]^T&-�L���`�4$f�F�d���P��0lB� �Z����7^u��k��b���03B<OZ�V#6��,q�Z��KA>$�C:]9���p�v[09]OZU�7��Pi�_Ͽ�e���g���I�庴s[O��2hMo���-E�	l:�:��ߕ�n�wd�yjE��f,��b��)�G�m��?���-���]�e��q�Ԅ������_`<Y�O�u9�*�֔�ZA��h1�	o�bx�2;�767D��/e��L�-h�G�O*�b�E�.#�[/�^$S$�I�p�5�����J"�>�،�.��yuyV�}$���ԴٌInh��\\J�ߩ2�P���/L�C1pH�l��;,I{_ž/�ͽ�y�%\���Tؾs�zFs��)��[?Q,@��}�]>Wt�.qn�8p��a?��s�b0�|H	�er�u&ɬ���aڎ>o���Lѱ���������;����~u�n�!��n�C�$�z�̩�L
��R�:yT%6�]-Ȯ�U[��{:M�fCF�J�L~��<�x�A(��f�n�%��^�������A�����R�����ѦF�sCMƹG-3��G#���YyX�Yv��g�>>^҇�e��K��B��W;��W�Y���1���#Du�*����2�3�5��Վ�B���l��D9f�SV�e�����
 ��<a�2��;;����gC��<��>Sc�������$�z�Z��L~�4��| ?F@����Ę��e�(��/K�3��Y�ǟ���ڻbGgQ���v����Ś|��N��G��9�_tۆ\�2S2�-F�mJ͡�d��y�q�$���K%�o���?Ά}�I � 7�{0�o�8�RF��Rw�4(G�#��+P:�+"�=ވ<���L��Kbt�n��B#@�j��@�6oBG<�V������s3T����Y�x�"0�ԏ���6�N+!�U�R&��0(锼�0��d$��9��64�qrO�l��6(܈;U�4���^ɿ�eДN������<~,(g��|ȥ�����%�̗�>��^-s�p�g���R;����9/ჸ��q���0�"�^r@wӻ������d>���,�ט�o�W��y+�6�m�'��:��ĭ����\s�R��(�z��#��*�o��|W�	 ����y9��v�`N�M��<�m/�uԇ���
!������#����[����dl���\g'���q�\��
R�F�w��;tW�Y�;�(K��:�͒P�%ĭH��wB�y"��ؕ-��~f������
��=���e��>6�����U�ǭ�f7��tؕ[��X�i�������&�Ű��X���Gɗ��g�44�6F��m��/��!�hhf%O��~\�x�4L�金3[	�])������P�(w_t\k���|Xv0��2�XI+�:��R4ڛNDF�����.VW������v3�I���j�љ�/�*��۬%�*9˒�	W��M���߸bkr4ᭆy0Fd�.^7`knT���؀=�8�vH�j���
��℥�U��M�=b�˒ho˘�;'(�\����K#��E���Y�C�X����b�q"�q�LH�;���)u�ql�m����eHz�eؤ~Y��D䜈�=|�&pX�C�	ھ�X��2��Oݭ�i ���Q��ab��߾�7������J����	sӲ�?lJ�U<\I)#�+��ó�s�-�!i�
MH��p�Z�����.Gi'W7����.�C-���Ùw� ���O8(f3zm�]�#ɿ��`2f�U"�p�?܄��S���x���<�ޗ���_	����Tm� �*��&�6�U�u���5�P��q�Ǥ䤘�N�bY��~Ĩ�S�X{��EU�S��0��Þ��v������Z��$�d�8p�ICw`]ny(��FtX�T~�u�\"��]ۺ�T�|辁�cp�[�ԉ�y��>��GVa�Jf���Q?����� �CndL�R|�1"=�g���z��`���Ogt�&^	��+n+��B/O��N{,�b�lX�G?�oZ@���N�ϲ�0�
M��X5ko��g�(OvE�Ν�A���'ҬH5�r�m� ?-�s�I}[�[�{ӭ�H�^F��ڵ��\p]��|�qx�N���-f��;!��1�"�ۤ�j���?V�qI�Y�Xm��o��O\�}�՝C� �l�!|�۵��j�v�����*a�Fpa���1h�xV+�xkf1Pu|�drk�����V2��Dҷ2&���8 M�vi��_�氈<�L���$@x��jN|e[�xR-P,�H��Pe5<ױ��U�\ͨ���R��$�k|?�����d����n�HX�ە��ПX?��&�ɩʃ�(^��Ҳ������rӧ;B)�3!+��yK#��v�c<�&8I��R{-#o뎬����<�p��*WV8@�1�؃D䰇�b��w	�+�����,b�K��%��ɣ�R���f��3;1 �@v	T�u���mN<J��(���ʱ�FM�n釢üf�x�ˀ����_P"2�)�`�(0�ԹREr1�
����ᰪ��7[�JYrcj)s�Z�7T�����&n��n�T�߅ỌS�F�hY�URr�.�7�҉M�ҞT�Oϕ"Ai9h2أ7�}���B���>ީ�1x2�}S�y��2�����x�� �Y�͕؍�b��G�PfW~����i���IH��l`��Js���*M��Y�hL�F�[�ьk�hb�Y�R�Ku\�������EzW�2�YXŭ���VI���¥��]��RX.Nq�Bu=��^�9a31����V�h������I'��"�C��zV��N�5��*j��4ڤ��ރN�:�PI�:��}Pt//�l9YN�Xq�5W(ed'�ԩ��4�n}��lN�Y�T*������/&�U�P�L��Y�"�ܛ�� Ǯ<;n��H�E���N!7�^����%��es=��4�s1bɖB�*����<�`o�g��hN�fB��v�"o�B�E�ˡ�dIG�9l�O ^a�+R27���`x�-�"�������'��>�T�S.���+#���G����i����Fk��|� !�ܣB���..��G� �o�	�z2�<'�h+?>��*F�?;�>0H�g�Pуx�v�k�^�>R{�)k�E��d�vY�g�G��'���7:!q�/Vw��}e�^XB��b�|��y��:��g�"���UVtd�4�����o����+��qrJ;m�?���w��m<Я�Ǩǳ^�Ln���.Q��D�TШ<~��;�D�ǲ��� ղ
VjE���O��|!��f&�&�.b��x� �y��u�.�o�}�:��*�<��	�s�U*ߚ9q�h�|�Q�\�&�#�}(G�[t�	9��p{V5�K{���Ĉy�@���Ȳ��`�j_ѦGu����� Eq]՚e�/�}��Cl�|.a�&;��{���aR�&���23L��&�^��N!;}�:�.��|ׄ�����N�z�wv�~���e���]Z
����h3X��1��o��C��ˎ��S��3�&%�2@Ph���Vc��(O7�?2Y�i��1��/�����<[�U�F�{ͽ��}BP����;�Pj�m'�M�l����O��$mU��ҕ�ϟ�� ݧ���ize7����Y�O��dBt�Oޟ�B�"+�O�u���/��ٽo(��wQ�&M�E�`��|U*�/�l�1���R����8�B�j�U�7|})�|߅�{�	I�p��}/�uv���lZ.vן@���q��we-�I��B�vQ[��B�s�Ǚ�a��]2�����'J�Q��G��"���K��e������$ x�2�EԕI4���01���6�E��0�W��wx-�3��d3����	���9\�r���3l߫y�9XĚ~����9�L�ʎ�D����ɕx/6�NP���K����v��g�o�J�@��q0������=��^�����[R����p��_D&�'�$�J&�^�i�<_�D\�������?�pF�ѻ�IK�s~�WW��B��]h�+��\i�fz��O:��*#kkk��9Z�����H��G��z(loB��g�b�> �bx6I��gWFʬ�E��]��[*�����!;�]���6�4B7����Y[�h��=��������>�dE�w��7���H9ǲ�D%��n��Y�Lmt�G���hĪM��b!	�U����{�^Fi��.y��뽦.G٪���j�hc����v���^�F�[nTBW�u��+�-��=_Y�i��;����V|neGUN�H�MPtsQ\	�]��}�)�0�<����F8:8�M���d��X�
w,H#�����|Ԝ*ȕ+�E}�"�U#��I�>غ=���rt�R�#��'���,�]��A�٤�7ʴ&������ �=⫱���	]��Ë�a�@�}g1�iF��Q�LasZc�w[Dj��F�/�k��3%7H�d��vӬ���d�O����ñ������bD���A2}�|�c_2s?MR{��,��3 Ťr��P�u��� ߔ�iQo��W8�j"v8DуX������IZ�9��%�6-�j��y��@��_@��l���!Y[}�3z���^�"yb�����PU���bv�~�fP��ԗ
����d<B�Q3��W^�ҳ��q���k>9��V՝*BR��Du��̚��=��w�����J���/��y}����䫎a��t;M����4���_�.=��5�Om:����t���
Z�qk�+c����#�礙6^�r�Y(��M�V�M�}=^dm��@F
6X��uw �\D��y��"�
)gC!o	��SjŻ�S�VOU:��$�&~1 �9QP&��r�`��Rg[���)��̛9#��"uR��1kӳ��Ƨ�p
QO`V��\r�A;g:���{1�z�ڸ~^Q�SD8g��y�+H��|5�I�.���x��c~P�M��r�̷(U�u߼,i��]����1Ն�E�	R��}	�r6����;b��N�'�;;��i�� ��8��㗬_B^��1��E�ZE���L�j����խ�Ѷ���\4�	Ԁ.'���P�ݱ�E��ұ�g$�]�:�}7��.��TS3�[�;��eɟ��,s0D�����4�wu{h�	c̦�1��95��!d\�N 
V1��c�Tt�ƳE��KV=�-q"�+G;S���Mi��Y���@^JJ6̅���۲ͲS/~�H`���*���!�?7P��TK�f�`�Z+��¯��iS�`���'���ӌ,TX��A�2�0�Ҍ]l3Ѿ����@4��9\�2��u���o^��^/)r��q�XL��f��g��'�,���?6�����,�	�����յ#�
����������ـQ�����SaAg��GnVU��ԝ 9���h���"4SI��.����㫑��+����vXO���d^�N�ʗ��ӿ_#+1n����Z(M::	Q��F#�9�3�����G?���gz�5��>a�iS�'�nsm]��s#�9Gd�o<�]��!끱��`!��xǓj�5q��C�6�8 [�)Wנ���G�(AmU�:�-��A�8�^Ek��쨢��%a~�-�Ӭ��;��^=[�҉r��1
v�!Ӣ>"AGI��t�_�*s�'��w������B3��>���ɬ`#}�d>70���2�኿VA6�~���io�9�a��r��y��u�7#�U_V��YW���X��%�����,F�h��(�E�Ǖ�ͼ�q�KB�K�~ݛ�``%�2��M�Jr�/1��j�cӫK�׵3Y-���۬�w���aMdj�Gky��/��=���:	L�&F�*���P
�8���B�z�j�"R&�'-5���ŏ���,ݙ��$���
�l��0Ї�Id��D`�p�w(�=�����ⱉ�~�6��S���MNJ]$�LtW�͈��o�[HE��GRS�wOr�"5@�X�`l�5MS�m��-D�$<��s��&�&���Ց�UN��p�M�dK�S��mҝ"����*��g_�( o	�E��^S�Ǎf׈r�ܾ��SO����z��K���4i�P��|�ks�z���+L��")�"'�����%���F��6ů��)�9EΈ
��J��D�GO���M8����ס���F4��f(�F��~�(h֠"����E)�p�+J9mn-�ϛ�=�t��`6A�^{w ��qj�$��7�!$̵��|ȅ� ��O�� �Զ}�}�xG��N�Sj���jL�N��@�j��7ag3
�4����e����5��o�"�!ٳb�T?_R�;�X�:w�^o p�1dZ`����f~]�O��A�u����u���{
0|��*3pk`��:l����uq���_��J� $���䔂!:$��˥�J0e�vx�ȹ�>ɟ2���1�,1Q�Z#�n5jRN��]B��Zq/��dD�_߹i���0��B��!��^���k�+���dgQjET����OwH�"�X�4��.�_���Z�R�&�]�,<�a���l��ME�w;���X�<g�����"����������+�ϻ@�ۻ����(ן�ka�{ɲ�Y�'�A��9���4$�s���-S*���(exNw���rGk3B2i��>����I�0���K'E��@��$D6�����<|�I��i�p�6����'g�[��$c��+-o7�a�0�񻏯�w���&X�W��I��iR�:/�E0��- �]�p�{�v>ZE9%��(�zǤ0���jH~���0���lQ!�G�Z��LK޺�|5 �1rĀ�mؚ�gl��޲٥"�P+���sUH�BX>
ewYO�n�����db��mR/qE��qEi�^�׭��V�+�4��+F�A�e��̹�u�T4�l���q�X�J΍�$Se�MQZ��hI�f$	y�T��w��M򍻯��@Q�FM�:����Ik�c9��S��rڤ��岀a�u����h�����L&$Ĳ�ς,\ڏ~S�V�c���.;&_�z�m��[�lH*�� _/T�O^$D�����/Dr�ec����	E��͸zf9��������V��;�v�u!{����ڹ|��+������.�B�%���
Ǘ8&����Rl�����DԲ&�ξ��x8��z�ŤV�>���G����� CP~)� ���s����5��E8N�,QvX�-[��u�l]C�E�2$��7>jo�#�]w��(�?�v>�@1͗�j~�A풇6B��r���>��G�-��Xn���ۀ�`;��`�@C��������8I��J��fBj���ݓ��I��LrU̵Z�T�X�	�7�i<(��R�~qTz��j�~�����q\B]�AC�Q�l�_��3�s�5��|���� �	!��8���u��,\Z����3^�6ͽ�CKC(�"Ċ��I���7�L�"cb�Ch�����7�R`�T��ԡn�US;兌Y8H���Kp_+��My;?�pmᝐlx�� mPဝ��V��uR�Vb#� K�>��
�U}Ud�YZ`?����$�]��F>9��3��fk�Ν�{���`Q ����|*@ ��3��*�8�D���V�v�I�����ЍQ����d���]r�(��.���+yD�'o��~��~�J�d,s��:mYY�FV�u��~�5LÉ�,�K趑ʽ5�,��\M3�v���5����Y
޶�d��{v��i�juf KM��O^6v���枞��8�t
�w�aM~c�Q��_����C������M�#��;���ޟ����P��
L�nR_�|���#�M瀯p�9��U���|�;^M��^�q���3�:F��0�)� C��H6%V&�V]m�ۏ�`��I���+��;$`Ч��e�z���>�hP1��}g��noH��8��uī|��Gc����޷��Ȓ����sᐋ���Ш�w��7�9�j�:w�},`ҨZ��P��i���
��������@&����5�r>�I�ZH�<`9_g47�Q5o��ɀ^����BW�O�Z	U|7�dh"�����r&[�'���N�����ڽ|<��Y@=c]������7� �� �n�0�
d��h}h���H��H笃y&���r�U���U7n�/��I���w��ӂKk��-DY�<Ȕ{\f�`�{�,ZN^A
��O�Sgr�Q�?¿��2^q�|Y����� -s`ݒ9�iD���6���s6�R���W�R�g6�u�,���F{�SP-<��ɮ#՘)٭m�����aBx^V���)L����( �R��m� N��a��ˊ.Z_�W�t��a��r��8�z��<vVX�Ey�8#��َ����}0��c���K���ч�@���>.^����D�܋�!WzW�MF
D:\JX�Y�Ni��V��[�UT3F��3X�/=�~��+������ �E�sg�h~��A�1���s���.���;�!@��[��P�S�� ~��e��Z;���!(�a�O��q��:�v���� ��d�����+&���e�r+w�-�@�Qaer�r�jDe�z�j�(s�!�����*��{����3�ۘ|�KbQ-�t35&�;��/����t;�es�ęg�s>x���N��1�͢��+���t �C�;ė��M�e�yˇ>%D +����u	!0B,:�嚥��̕��Ֆ�[���΀��O�1�/7�!@3<�BK�����j��A�	'�W����y����"By1u�X��%ֵ�変	��'�?2���r��5M57`�m57�)�W�b�k8�Q*���<ʤq;�V�;ڍ3D��Rd�7�`=�!?HD-�<<R�k��hRV�LWV1wPhLN�Q�>�(�rl� �t�8�&���!<o������M�B��X.�%�SDe$6])��bڟ��ۊ�|��ksQ����CuY�-�m����Onz��<Qȭ�C����oa�i��$�yӳϱiV� Q�3����o
vƍ8��I�-&A�����
H��b�/ߢ�"6,ccm6�?�M�_:��iLX���ɹ�湆bYP��D�|E^�;�wY�̈��\��ޅ�g�)-�3j���a" �
Ra�:��a_�h_��D�/)�U�+I�*>T���#lG%�P��;���l>r��i��u���\bڞq�b/򊢥��̓9��u�K��"+�?�jh,�ͯ�@��aMh��SM{�<�D��8.x��wXĀ��}�= �X���A�)���j���y.=D�X�,<��4��s.æۭ��ρ+TL�0�챵Cle>6�[�O�Q�f�F�%!Z�mb����7nj���+�<�����1�����d�V��I:�.���|8Um��w�F����ef9 U>��,l�E��x29���:�,�;��+b6�3l2Ť�?V��LZ�fE�`��sz��Z����U�H��*mk�>��"��Q���v(��05͈]x��e����+��@�=[Rih�K~����C۞��]p�#�������f�|ibb[� lRz|W ޥ��h9F_�ỶT�[c�l�������<�s|��6Z�-��m�}F-���q��-2��C��iH+~-T;�F����q��v�h>��u�F���#�'�K4����� ���yH7��C�Tؖ�X�&c��6[?~O1��ط��Ԣ�}��������_�����*���t�E�����ť)77��L=j3D����n���h�V��QΉQޓ�kmo8�f�fA�lJ��s�"��l{(�c�� )t/����Z�������C1���>�Q�
{��i�@�{<G})�G�K�ӆ�$b�7�ŝevzd�ftq�ٹ^+�����ܿi?\d��p����'�{�c<���<��S$�z�������0���R)����wx ��Z�|�_� �e��N%��`˿���2��2�8`�"j$I)����5���_��h�w���
ސ�)�C���7���R����CU�<z��H��!���kQ_�%�0	��� o^�@�M�o��ڧ�H�!s����nѤ�|�C��i
��!� 
���IL�294Q�) ���o�`.��z�����y�=C��\:��� �T�bhI�E��.���3O�����{d>y�>�nc,�"�!zA q���=�"j�Ȳ3_þV�*tA�����k
��ձ���Y�gb#0�M%���2_�k�6��gK��2�LDp5�P�:"?���!�[�LmP�QY䛳��-�C�$�ԧ���|cz���9p蠋��}N��ia��-�,_Z�N����q�S4%��Rt�������옧���ӟ]玥�`�����8u/��zĤs���t�������o�"o@S�HHe(V���J#��/r�M=�o�
���:r���ń�f؋#!+�����������`���!�I�t��9�nK�5�4��Z���Lh���r��j����B@bO>�������73f���Q�:�Yû%6���z�ɬ�&�D1z��-�F���I�]��Ú�ޱ��rx�剄O�{'=}?�ma�U��M�O'���7�5��0�;��U�z�"��9�G��\�C��X+4Cs���S���iT��0�����8B �Y�)N�X{��/$׉\�Y7�?�}�	��ɉ`UQ��x�[˺���7�N�5������z%b��~ȿ�g�)f"[�~g�|��yk��v �K�^s+�+[5k��GI���Wt\�r
^�]qVl�F���쳨M��'c�D�e8�}�@����=���	��Q{�=F�_��4E�[3�vO���ߓq���+�'��R|ԵY�A�k�<,4�Y>Ժڪ�nPo�q�s!P]�
x��W��O�2��Fݣ��*��Bv�_�B��+2UlY�;O�䧹���b�����O̪��B4޵Ը�n�v�Y$=L��'[4L��ǒ�2��G|KEO�.Q�S�F�gFY�#b,DL2�d��|��Q��DSat�У����tut���u7�v�`�禵V�J��-|c����a��:��IҮ%�`ZL�E���a�w������1<�3ƒ_Z���HX-����̻O�kb~v��\=���>��?%IDT|&��W�'�}Or��@�|5�Pҷ@O.�R���c�d�w!M�'��Pusn����D�୒(��y ��߂�JX�� ��yʃL�贄쫁\�
����e��H��-�\�zI\�,*y�L~	Z��<:�Ǫ�o��B�`.u�XJgt����?��̘���o�u#c� α,:�p2`ǃu��I�cB|�֙�a,Fl�3��w�%Y(����,���ʝV��6~�)e����)�Me�T���m��[}�i>�Pq�aOr%ڔfo{T��!C�e�)���F޶�����4�LU��G�/e��C��n{F�86i��#���@0m���e͏jc.���1������@���̟���<��o��C7s�TK`�K�wK�|m�Je�8����6��Vˤ|���ۼ�]��Y7����� '�����1���8��]�m��5;�d�����G��]����R�r%���v�ǧ<�\b<��/X2S�P��.պ7s��ȅI�%�۳rbE��w$�ÊX �q�`�a9*��Э"g5���p��bkz�P�?6<�6����тܶ_��ޚ�G��(4~����n�`�$0���N���*ǲJ<�B,5�?/�l�Y3���V�wF[�Uu�i8nO�<�ҙ9��i�̫��1	?=�2�"h�e9��m�F�h�]��е�;�-�,mt�Q���7�o�{�j�
*L���>Y� ���<�����w8��3ܴ�`�ծ!�0X���*�a|�j�2$S}Y
��ؒ��Ǜ�V��K\�MտomU�yJ^|%7�Z����O��JF���L�/^�D�;��[���U��^@+xI��:, ËN��v�|�����5
-Ir_��e���B��sS�:!Z�q�&NR���[��-S�sf�Ij��dW��3�ݶ�P�_��0)I�.��2!`�V�5�E9�Bgz z�}%��/�{o颋�h��ټ4��� �L*���	���bf7ڒQ���=�{U@�>G؞��h�ݑ¼��!��{�3���o�����x�5	Us|0�܊A3IL�w#��C����	o�|����'ٜ�Z�ǂ���è��=��LW,��}6���6�[+� "S���*cW%k0oK�b���~�JR��l�ۗ�b��e�,���g�J8]LT�b�ҫr����8��d;��K��\�9���+K����(��{�I���}Aq<A.��|mw��.Yf�z��9���F���t��n�]c1����7�b�)-�⑥��U$�@��x��I�=m#������~U�7I1/Ӏ
|HSO=�d����v�����m�(�ݟK�t��0�v:Ɯ�n¿��G���p�R��?�B���rS>E0Zk*O5v$�DѮ*r,3լ5��ԏ	?��8S*�{�(���ɽ�.�Z���Y��9�C���O�
V�� YB▯:�h�q��Z�q�R���	Zb�"�$�M�#K�����[�M���z��vf�f�~��*=f��Ps�f�����Jc-(�����U�E0�,u'�/	��q�O��Ǯi�}��ͣ�ι|�F�i�3����@v�C8P������ߴ��zQ!�6�!���V*	��5~}��\�4�8���{����	����tC�$-���[+9����Hn�hR� ����O�&�p�a$�%K����
�hʃ�`��JtSL6-5�3�(�>���pJ�/I�:�9}�	��Q�IV�k�u�p��x���Q&�#���ѕz��j�ݤ�������l#�[�e�(��}���aɸ��w%��7I@%����0�i |ǫm���p"N~�mwh�k���7��	�?6�m8!\�k[褅A?��=��2���URBq7(�2�y�Wמ��l�Oc��w���t�$�8��џ�U��b�<�;�k��Pr��(���6�a|+�"{ԔU��?6�dKΌ@�-��h�?�����!n�]"���8+�K���\���H�����&�d��*�P�7k�~�����e���Nb���ƙ:c�mH	ooxl'�ف�9��;���0ZB�=��@�����'��]"���~��|0N���̨c1L���(��OK�wnK�c�)���
��I�yT����//T�`�*�"����c% D�+,�?�����D4��S��e��& !���������p���8�օ�>���9Z���iY��W����=�4m��$��B�.uC��ꙟՈY'�����Z���Ֆ]����+J~ɟ��D'��Eg(����9������c�"亨)���X>4;��؃'�B�UeZg�x���$d��{j�|�
��K�nEW@�ZI��3#o���[�l忍��M	�2��>
 ���d��A0����9s(Ls��G�)�]`3��>�$Ya�`G�]�����ш���Om��qV{Y<�Xg�
�TX������Ј��ͥ-�H��*�?B�Υ��>Y<��H�Ք�)*���?w��)����!�-�	GW��0�c�i�b�PY���y�����٘.X�EaHe�J1KpcQ[�u�3�� ҟ����Ȍ���,E�2�U(��Ix���$�o��\�Q7��g����NSP�+K�(y�-N�'��M0�j�^*ƻYL8X�4��}u��K�a=��߀V)��a�ţ�(;-%dc�USnߖ����k��{G^��q9���fq{��Y�j�X �6�1$˖�ΡiR�>In��}�@60��V_�9�3�k��)����"�t����7s3� �BJ��0|ñ$v��*�ݠ�("��I���3+8�;ϛ�=�&Yw�`�SӼc��������g��gO��ة����vx
�X����2C3{cہN6x���$�]�����U���5��r�rΜ�$�[�@Hb�P�j3��l���L8v�F2t������+�����mړ�:W��3�Z��\�憲�����gu��yBz)M�$D���7�)o��A{�ʍa�l��P�eqM�B=�Z�#K8w��O�*�ǈ�;�%/�]%�S����*�%��-b�bU�R�eM?ݹJ{K)�g.f��$YH?���<Ћ���x;+�<�����y�m6:ؘ���z�$c-���W��S��lSq��&�7���!ܓ���[�VS����tAcqzԇ��__���(�>&/o����x��v9ȉ��l+f<�����?�Ut���A� l���y��6��S�ٗ2/�8�;�-��H"~4�L6%H9�4A.�<0Iũe*y}��I��|pa���9H����\���04T�x�or|���:�	���]߱������\������efrv�!����jEz*�  !��\&�����wi�i������g<G���	��$uJ�]���-���BS����}CE�c��T.cv?M;�X,M�V�	��
����Â��!yc��!�:%C�s��1>S�J���D���;vrQ���.�I�H�H�y����R�6�.|�8��)�׮[�zy+ӗZ#�ޜGu�A�ʷ���)�!/�x;|�6�{�p�i��^m��ԇ�����7�������$���4ޛ��R�.�����p>'��Z�&zߨ;�t���;X��2�s���]���A��X��+�537JC&�և3�3&���d�OtG�Ǻ�1�wl.ઉ���M�޷�F�a6�!�ki�;��y;����<,�נ4��>d�M+ل7��	�y��R����9l�,���q���5�W�oP�!\��c"}�x���ԃM��*w�~m9�o>�����i �s�!�X��_da<��>3J����AbJ�A�ٔ�%Tû�@�Gȓ�@��H����A���3'\����ϮO��6fh.����`�*��uJ�1h1�ݔ���?ݙ�������<�4qG֌՜nۼ�fâ=�,��	t���g�>�´כx5�[ 3��Aԋ�{f�e-��F��h�܍�����>�E,Cs�c�0��y�#q�9�hl4?�Z���t_�&���-�v
���-�:\��E5��S�3��#���|��	rO��Q?$�֘�v�#��ki�0�d���e�0ޢy]!��� 5�l��Q�f���V���u�TK����:�,Q��i���"{�~���)�Wy1����b���u�z�ف#<%�B�6>���6Q�vϢ����eq��P��H�������5���½�[�)V��!��M�E��ga�����BfQ[qc�6͞�p��x�HƜN����tr�ca�	9{���|V�=#��G�K���s=��\��m�N��O�T2�'��h.��[��4l.�ě!��7�O�\K�q�EZ�29�Qy�8��|�y�÷�A�I��̀p�m��׋ՅR�����Ai'�O����x�%

m�Q~
�>=��R����ɿ9ɷ<d�i((�p�X���co޲��#�'�������.<�Y��de���T����,d�)�*�l���>�+K�rPy15m�o�`����+MZ8)��E_�F��/TO��ݖU��ZKQ���1��R��FO�$��έ�ke�؛�`��
�f�e�D�ީ��;����l�wV{f�rޤ�t�ʻ���Ӳ �J.��P}�PR�BWӪ��%�v���'W�L���G��V�<z#���)���D�ɶ-��(��ٗ�S!T/#Fz���ŋ�d�׏�����^���+���bRp�����^���%���+�
Tn�����ĥ' M�:*�i�I��X_��b�/��4���~*d.�7��¯�A���T�kq�c弴��0`��B�ŗBpC�v�L;���*���:�O�JH�WP�����E2j��� �Wh����}֑�AU@�]ى����8&�#)Rfvq���Mczv%���r1�M���r/�x�o�W;lH�FfA+@S0�o�h��,ӣÆ�7��:+����u|�*b�<T�
ҋ��w�r����`!8p:�(�9��hqXI�B\��El�Cn�db$-�TX��g5`[�(��_>�(H&�4o-ߪZm8�{ck7����n�t惥y}Q�v�f��2�{�sDT��>�QrYy tү���:8�7y$Q�����S�/���WUfʍ��S	�S�7�qk��h�%3P�Q�ɺ�M�UqƘԛ7�b�*_}[C�AF{�4OE>b OKG�~�$2n����T�"*K��A36�U�ٍ��[�&5����a����T5^ ��MI��'^a�М1�
i͓�֣���#W�m��9V������E�
��]�l��"���3$[��V:_�;IX�?����YInN�=����W����$C�#@uo(K�ٛ��j���X�䳁���n6�^��:�g������
 �[[��f����v	�p��"�Jh�%��J����E�iVzT*��z��.j6,$��'�����:/�b�O���5�̅5���C�[t������#`R��M���i�)gT�6����B��덩��,ɠ~�� �B{	��*$he�!�3�}K�t�N�%�=Jm�~��@��!�S�O�����!��i�ɀ��U�HU����ؑ�Ś�D�q1�����P<�k�ud Hg�<�q��]Ē�?�"0��*�f�h�������F�z��3���I`��<�՝������3I��O��&[i7��@�`�*p,��8ǟ�H��/n�6�tۦk��u-q������ێ?�aw~����xg��3ʶ㨫ml��ʅ�o����P[~>K
��P$�� �/ÑJK˗����}�x����}/o�֏�`F�&��?\,��F~�_���Z�G�P*k��4�	YU��`��b�$�P3��7PYo�m��j ���5ԭ����y���/\͝�]:_���O ��K' QĄ�=7�q/p�zn��8hӞ���Tx\�H80SvJ�S��	a��s*=�=Ѷ*�u���&������!pVk��5� e���|"+`o����`�n/�J��X�TN!+��R��V�����%�+�n�J�	�����Q8|��C �]x+��έ �WϚ��`�>����Q~�PEU�Tw�"�B���MHd������=[�0�|��ζ�AV�8�=Dq��.�����F�w���4��D�j_��u�%Ԅ��<��]E�~�����_��sҫ[]��?��Cb�Q�m����<Ux�v����xQ���v5�-|�y��!�{'�
��yi?HEg����!P<�(�>���aUh�k$�S\}Ax��'�;h�p㛜�LK�+�#MUSc>���^����@�eH �2kO粦�I5\i�x���w쮓�B8�!�"LAw�G�q�:�g����v��#�=��f���p�k�����y��@XEXX��$��H���FL�^VO"�3p��{%���%w����D�e�����+j����FC�%���!�1�_�2[�r���@��ȏ�O�`�`l��Nk��9*SV�-�������!!����~�\�z�N�C��V�Du�/�:��,z�H������e�S6ٓ^i@�y8q(��:��M7��K�8��5�/��(m�c5g1�XF�"}��=C� v��\׎�ARҋ����_;�M�S��EԽ���z.��9��L�Չ�[��?�_���Y��<���ܡ@J��|����b�q1�
Mn�qѦ�I�O��� g�H�r�K��{GEOj�����h�Ѐ�ʰ�f	��V��� ?(�/���ۊ�kZˉf�c�mۖ�9l`��.}♀#��賗�1�m�+u����e����'�Z�T��C��z
s2B�R�|3�ה�[���t� �צ������ݮ��B8t������>`R��u7>d�D�#N�� �!����f�!ʨ�Ų�	B{smq
Η��o1n���-�\v�]�au�����ޘ��Nچ�ӎ?��H��z�up{�������p2�fB=�� �PZz}޶3�X�o�2�nu�)^�_�/z��Q76s\ޓ�h�N�mL����a���m��"�Ϻ��t��vHE�V@��UCE�=�Y�8Li+�����W�t��|Y�O����u�&�J
�S�����i�uO�Gj�yDR|�܊����߯�ƅ�h�w� ���*]����f��2b�s�EE�ZM�ɾ,�*�&��-��g	��G5��3eW���� �xR ���<�$0\���X�l�O�h�X��t}�f�'���c+�{�������*^�5�:D�q7@����ȵF�d�y"e����,5|r����!�~��"��\hP�*pN�A�m<g��f�%t��y�=B뻤��������zlJV�����z�T�4�f���"�[XT��+;BEA��k�1��Y�exl#%+i�����vDҐ�����zEW5'E��	���\���y���s�H٠]-/��lH�.&��~��	3�������o�0�A���e�)(�	�0����C��-^� r6:^⻃7��m�zd��ɡ��̄�6��Ui�?���ơ�'��8k,�Y��q��9:�Ct�X@��xfM��S=���I�� �Õd֔����fe�z=S>�*=�*&�k�\X�/����5��`�|��S�o:��0h�P� ���\A�8��'�_@O�'��EI�pѿc�p dX��Ҽ i��]�<�P�_	���ۼմ�F�.�K�(�Syi�L̀�3J�Q|�M<d�u���
Kl����� ��L��fv�%à������^��<�P;�(�u�����G��+'��{��.��t���CEO��ɬ"W�9˼}p[�O���"�fR@!݄#�x�)��F��5K:�O:Q�<���A^�{����E�����#ߣ���`�� E�#��;�ޠ��ȔET�(MB ����KuJCD�=y�b���!0��s����ĸ��0�D|`u�=���|�LX䉍�~�}�l?��4K(�4X7
w����.ۯ��P���>����?�md��y��%���6nvĭ�1	���	4����$R�ܙ�w�A&��X�s����2&2�)��
P��L��Ioa%��}p�䉇v��P���"��ˡi�[���6ܮ��{�9S�$��VV���}��ބJ�<�_�c`��������VJ���sE�Q,���-�`�M_7	#�K��_�ː��a����BKL�
ȶ�%}�&��&�	!�0��g���{(�����N�Ļ-�W�e��S��* �wz��{w�*#,�V�4�Y^�sԟ?�D@׊)��G\�HDǮ�c��7/@�E��A�F�6RQ�9c��$^ ��<�� Piζ Hhu2N�aE��Ժ����+�)ꈗ�}̝w��{bٯ<#(ض��~�&�ՓP)��d(�Nъ>�H �x��ϥM�N\"�����W�.�f�\g�6�ᛶ
i
�}GԦ�uCqu�/}�&��Vi<OL�KMj��,=�_A���~m��U[�ݳS�K�_xoL�ڨ.k2Qٴ��*sP4`Q�+�ciG���ë	�Ps�a��#�ξ6���EA�5��q�&x�C�|��x�;�D�
���c;���F�d�� (0�{{Pv�#�����$��G���G�9�챜0"X��9�(&�Y��ď�?Z� ���i9Ιm��1I��&]c2x ŉ�k���%&f������T@�c�Omr��%Rx���;_)c��G`+�f]n��$���ѩ��m+]�%���a�e�u�c :���R�-�,��8�K�:�A�|�V��d
(���Lo��C�,�`LvsC�}�	�QsԶIo�Xb�E]�_�.�����u�S?q�8��j��WD��wqU��nL��Ѹ�0�%%	�n�#���o��}\/�y���s�fÑ���B0t^G��Ҋ�T��:���Ϯ���f�:���@�����[N�~��l4㈏_�V��:����|�(��`/��`�c��N>.[jw�����+9{*h������ɪ*>.Z2W@\rl��CHN��寉8qP{�����L'��N϶�z�aRP���",�-Mr.I\j,��;��o�������H���bp�j�;L�U$�L��6Hh2����V�vT��B(I����c��(��u��*X#�\��s"��m�E��r��t�d�zZ���$���9	l��7X��Н��z�:V6\�Ͽ���{l�
�x���	TM����ĺ���Ƞ���j���){�`�4�5�w�"��x��?f�g��O����1�|���*�i(��r�U�[���M;��~C�P&����>��<J�z��3`��q���a���S_�AiÓ�'�� r��㼟$��	�h�X�hxy��˳3~]gd���0�� E��%.)a�R� �U[��8s��J���2��(�5�ĊZBA���}�Ѷ��~�'�q�,�ь�~E�m��_|j���΃�#^�dH;@�=�L!���'D	����4!&mQ�����NI���Rf�ctk��Yb�./�賐Vo�Эu_�~��ݡ�@ְ�� �I]tp"�7mH$~ao`��@N�!>Z:�0g/)F��xB,�v]�T=%I�J��vMP�֪F�m����:��m�f>��-��%E�
�Y1�Ť�R���"��&y�̸�VWr0)�ey��gV��@kP�M���`��%dm��5k�r���3���!՛7�f�����t���s;p4����N�|^�7J�5`cP�b�����b+��B�*��L��)R�c֙-��l��hJ��A����@�[�{s],�tN(�w����Hp�2C2���:�X��H?�pF�b�ρ~p�.R�8�}X�GK��A�N�;���Tf������pW���f�����