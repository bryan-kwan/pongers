��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)��<�=�!�r�eU{���B�{�����zm=�����@���`�?vj\��h�0�$�j��W�ɏ���1�k�\�H9�(u(`ف��^�?�;���h0��_��?�!���<��7}�&�G��8��zt<T��XgnŁ�	��on�-b��cj���*@��/	�]��{>>��T�Gz2�ڄ�Z�<���>Fx����a���Ӯ�$�����]�V�Y�I�#��۱���VYSb2�~��\3��E���
��< �X4�x4�P/�e��I\Oɯ�(L�/��]��ϩ��C�>whAEy+D*p��\�~!�3���c1y�K7����"��?�w�n����4��A���哖�_و�Վ��
��`Bt?:�E�q�x%m	��}�FC�)/��SՋg9H�ϗ�z-�t����2�je��@��Ż�C>�x���'�8%B�'�mŉP�'�]M���܌(���^%[y�	JY��*Ҟ���XHF�b^�!���?�y�c��VC8zTK�//k�&��yL��b�!}�ID�ϗ�������ɳ4��#�:��͸��0	^bPB${���4T)Z}+3�f2f�Fy���Ȅ�2C�6�?[yVَ;,ˀ'k�?9F���ొ4?'��3����8N����g���Aiu日&nsP(#J?��n�a��zoj�!⯢yv9���_�\���5?x��Vw"F��,���?����Q>��bIl�H�<e����pv!:{f�9D#M-)��]Olw�
�����HW��R�I�(���ȏW`�%!?	��B��'�uʱlP)�7b��@\�R����������}v|5�&,�f��}&�� .��(�d�
����9
���}��;`@�#|�>uWL�M/U�`���̶r���k4Ty�Η = Y�=�_�>C�u���a��Y�%X_���q��X��¸H̫y4�����M��9o�e?��~}Z�PY~N�5[�����M˹�T�?T%�x��~4s3�b�?���q�q�ܨ�@���t��RWMJZE_X9'�B.�56��M��ϹI��N�o�D}� 'P*�T�x&?�X]��u(!�����։4Xӏ��Č �c7�{{�u`�D@�����阐�^#z�Ѷv�e⏚�,�e=�*Z���/�щ���`\�2-7r#��^�w3���y����v+�"_�MM��Bd+�i�<�hI