��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�����Ղ�vzl�br�6[y��'2�\s�2�H>�y^��2
�²���b4%����g����B!cm;k�w�;�ӯ��cedO[�8���C��B\�l5�â
����Q�>eF���|6�%��]9gA��Vs=x��pJ� @��B<F�c��Dr8�[Z'Ag�F�=��{�ߑ�5��+l�/�_��;7O�ǫ�)b�Q��[kCy��䶿���~˂J�	|:{n*��ϵ΁����G�wO�G��
Y�~A(��]����s��\�u�i[�V����},��WXy�Vf Ue}^NS��525-z^�Ѥ����mw�S;$�ݝ�1|� %�}/+q�qY��DWpd�z�b����g����py-]�@�L�y`��g�L�OkP�L!����x�f���d.����츟��O�^P��R[5
���~�W��Ev�r�#�b�D����y�Nc9h��}��_lXS�h���i�ػ[��^�N�����}8�v�5��h0&���
b6�έ�:_��&�If��*����A�oq�P�On�B���1���	�hT��*o�φ��Fw��ܕ�t����-i'Պ�kEd"E��̴���)��9E�_ t,LӰe$�������Y�����Ҧ(?H�\����~��j��c��u@~�Ǐ���-w+��YcX�����������jF)-�M!���B�a�G'!�$��Qɻ,�!��M���N;U ��(v��%2\��ܱ�Jij(�� ���J:���$?��ݣ��
���c[���Tʍ�N�hQ��\T��D���TӁp�;��i��&�<Q��s�l�S+I����w=��`]��pae?��M�0�m�`D7_���G�}�p��]��=��m?^8P2�9�ԥ�x�&x�pH�I��3
��>w���lPI(��L�*�盠#�m���H��]�Lf|+c#��	�`�V]E�{�tt:�[�H����
yp��r7G�*<����DW��z=��`�9������<��}+jZ�G�ߘ��ԗ�v�|���&a����3����������^/�ۂ���ٲ������㙋����׉�q���?<����=�e��>��0��u?�����W�֙D��V���� �e��xX�f��B�p^zQN_o5~���������+AMܣ����z��2��a��F%���Z}��-cf-��e���4��\>a�Y}w.3%9˗/����Q��G�=V�%^�����o�k�/��d�j�og?�*Г�����ǅ���:#Oqf����2v�Z��q�@�=��}��6�K݊�q�&���o�,��iR*�z�3׆k���.pMt���u�oP9���z/բ��p����o8��k���Aٽ����z���\�|��U\A�`��њd q�������_b�N�N9EKZ7�>D�x�.�������9a�̜�ER���l�3�5z�~g���Z���95��)(��ܘ�-7�l�t4;;m��P�?�1��8WI��#�\iv4�h��j�����)e�D�U`�rSm�iKh�%h+�\T��Si�B~Y�N�|ãZ���7eZ3�cы ߓ-&��X����c�3�|Cn�X�8v�;mDW�ʗ����x�q�͆���I���+g���;i��`N��qx4�6�l�2!ZcnS
p�&�J�97>߶r< ?�����Ma��W/( #/ųM"t�m�C ��n;�\!�e�š���%��3��~)1_)�[؟J~�m�3L!tN�VJ�1|�H�eBf;V��-駰P����%����3�)|��Ц�ʦU��N�:���t(Zx���5��Qbhܙ(�@��� ��U:E���s�a���lm��ꐕ��FXu��u��F�-���'��e����O����S�}r��L��STjyq�&����G��qcj�o,��7�|�L<� ��Nr"z�r�qR�YD2��/V�F�+�ܗd)����#�	�^p��[�����id��ccb<*f�_�^;j�}�M#�Q*�i]��ՑQ6��t��<�ݨ�96r:cg3����|�Y� NbM{��d���X�i�h����2[�P0~ȥi�)���6�|J@�"�q w����(`���{�D�B��ف��P�2���Ț�b�ĥ=Gz�?ъ~x��|�0�D�^�#��ݨ��8@A�Bdc�x��'�E���Z�u�f`~P���,��ɯ�PG$�܉��2��i�$�jڎ�Cu��^׬�HG։�X"ʐn�9���W�4�, �n&�^^�#�א�_R�X�8��X/�u�c
i���; �}{%�%�c*ɓ�YC�s*9�.�C�'�-N,M�g��"&��8�?�`��P���[?�|�(�
F6��au,�� R���.�{WE=�%�A+����q@Ȩ�[FA-�40�����v}�lo/kl<W��â��F��6O�עE�ӽ�Ox��%dP���ug��S��T9�\��B�$P!Ƃ���:�����ts�T�%�����}@٬�pZ�����j��1;N�	C��9��Խ~Dg6>Hk���{W��� ,��'i<�`�G�'�M��g-��6�L�|c-�p�F������3�?3�Ώ'�;P� �s�h��N.�"k@��� �7�C?g)���Ė�LN��c�#����"��-U;V�k;��/��u��!�B���Gԧ�1�L�ac�QC�4���=�(��ֈ�Roc����^�v�"��1�u����g�eHt�"'�5=�拞HNH���{�5�[G�t̸C��9b���t��o]Q��m��t#O�ô��S�:��R�ӽ�<�Mc$?�d	�Q��㱋��u�F�B=�-�e�����"^G@��	�Z�#N8��0�V�K�忌�O!XJG`e�!fL�#��L�wͰ0�7�!gt'�1�+ZϤ�%$�-AU�\8]'��Hav|9�k(=���W�VO�کƣ'$�/�v���)�������N��"aڮ��_��N�p'��� ��D�����/ux3x�׾�e�J�[hH����"�a�N�O�����$'+��_�ER~ιN���'��ܻ��Q0�w��;���?�0C�0�0.{1��s�Z3M�>I�^q�fdO,��r��Z���b��A��o��]�`m��@X�/\OU@b:s�Gm��>�A4C�9�o �IQ%z2FrY�A� jjQ۔ʜwe�`�y�s~�}�<~QFc�L�͎�Ҷ2]�y2
���'MP�Tѽ�/|	=mv�&���0��k�HX��ɇe���'��]!�Yd��)$kP3.��G�V�@(������njB6$D�M)#f�ƃ�L�N�e��i;w��i�r@����"X���H�ˤ)��:���ʯQ�Jgu^[<���%���l���F�YN��$na���o��K^��g���-�O
�2廙��aO	A����]?��l����,��]$�E�����7jm;&bd˞=K}��2v`['Y��A���9W��D��Z�$�Ȩb��8}gz�z����ӛ#�2��;k�\�Ӷ(.��ߏ������ˠ�簴$w�|�¬����M��`����Z[�����F����^�"-ˣ�m�H>4)���a}��������!����;<�
r�c�}��r~a.B���y߲�ݯ�|��4v){�M�K4v��%5l�f�&}Ԙ����q{u��y��i++��J8��.�]�c��:c�����������n�{�)���UZ�9L�I��6�#�8[j��0N���_��[ua�����߲�9e�p7tg��s\Z�f��"�0ڇ�^���P}�\!��w�։�Vʀ��Y���eOf=
eF��@��p����Ͽ,E�bS��Fx��6�ͼ�>Q��c�K�Σ�p���-������N�r
�D��(0�zٽ�j�o y~�i8ĵnH�#�#�p�#9ާ��N0�޺5�j��{�^h�Ch�:�u{c(���a؉�xT�M����]u���ҤRm��)6sGIq`�k	$*lj���~Ո��qsb���Pm
%Л��cB��T�v����H�~��`J鷅*t�8�+�t��riKi�1f���CA�h y��6�P!�/&�[����r,��O�N<5�G�@��'������J��F�l�%ʨQ���dQ�nx~�h������1*�~��¢`���)E, 6�7�x�%Lޔ��d&���x~�� mO�C�FI��;�l62+,�2'������Ҕ����<HM+E��dX�*�4>_'aK����c|�^�km���H��	�
��}`�ÚJ�����}�|����mR�ꪹ�+� �p�8�?��	b�I��JU�Ѫ�<�qVZ�Ɂ�ʏ���K0��F�'��&���v%eY��=��cIl�Wq�P�v�@�+�ڞ��C U�T�qa���5{Y�L�3��(�Y�z��
Mf�a��t$�� ��#7_Vk�x�S�	�F����b]�g!������ �~��%��.�A�<	��Jd}����N؄Ȇ�1�Cg�I�xV��Wo��\x0��4_�R̭ڢ�Ͽ9�È�(��2,u⿏\�
v����0�����~[��JE�P�{��d5�5��~�R�h���0d��ɿ�����ԴE����,�?�"��|�''S�U��:�b^M���P�T�[-n�*��A&�?�s坪���%H��IŶ�����e35UnJW��WR%-�Df��y�-��Ԋ��_� ۜ�o_P6�aKq���=�T��WST�{�����Cl����c?����pz�R�8��E �A@�i��Q�z/�x^tj�l���͸d�QS�&!����Cd(�r4:�&`���WTS�L ���Q�0��sdղ�.X�ix�̖Qբ_�=;Գm��5�R��t�Z��Vv��C�ݘ�ni�jxp�G��F��7�"�B�-�
�ҙ	!��ta��)�%�@� ]��\9�%��bXx�L^󰿞$�I�ڗwR����'�;�`h��S��г��O��Y���Z��S�Dn��X�)���Uy@��-N��h8�L(ķ��4M���[PT�R��������A|F}	��=�z�9b�'qQl���i�Z��O��p���\�:���=��a���k4�Lġ�����D��� |���"r���<M��涯C�2(>����UPf�Y����� ^2o;5I*`#AƑ)|�[��`�h���.���ou�rI?�Fe�ƥ��9]T�!��zВ];F��to&�k�J�x�Sɕyg��g��9�"*�8&N���NV�+�IV"�THy#x��|x=L-��U�R�� �>'�M>�b\S_h��d[؅��	�f���^��D��rX���u�5�fFp<2���3���y��5>߶�6�
�U{� ����(ꤝI��T��]��/����j�4���RpF�{?fs���92|�l�Y#-�Z��5����$�ұiv�<�#�"<y�&�#��0x�ԎK�۳t
�'c�5��[2:���Y����q�87�	���9Z���E��]���|�o���ܳ��M����_���;��,C�x����#��5ҿd��s+��H��$�Qx���|pB?�.�%���b6���+C�"�4-�"�.1�*�K#���d�x�q\{Ү�Jt�޲���ovѐ��p�7�X�L����N����r�1�eS~B��
ȴ�J~n� ���'x���o#����G���	,#(|�S~x�0��e��Ҩ��46�j�p M�4 �c��%F�C2G�9��oE
�>n�Yr����g�qfVB��Vw��VXt�`�궠�Y�6�آ���|v�6�~]��ʥ��Q��ט��r3�$Xl�G������_ɛ�/Ë�� P���ܥg/�t���^�6��^zAQ,('Qmݵ2�z��)A��c���*]�7y�Ck���3Gk�˾2��/���h��{8���Ջ[����QΠ�~(����_W�u1�R��;���8+D&@6+N�k}
�g�Zv�� ul5.R(�E�rC��R�@Xz�Z��;�0c�J��I>��G����ۘ]9&���ȁGmf|�$;�a���h26��D�'#�oWS��5���>��ϲ̕<�w�����~�����1`O��#��0�&�j�똭73�n���岌�O*���9�9�>]�/��|��A�z(l3�k����<�F`>Uf��!-���-z�����쾁�{)�jE|�J劣xB�wS��ahg�x�r���O;�4�h�C�&�ż����\s7�LJXa���Y��S삵ظ��nG�H��'����Z��caݴhM6���*-�o՗������9A^j2>Z�q�}MQ��~%��#�-�rY�xXҳ� ��j�;T��4�Njv;��w�F��q�d�K���M���4�P�㈘i�����X��lk�F�!;�(	԰� 9F��pOWB���	���Qf���� '��u�&
]$��B�o��GK��Kŀj��m��
G5��>�������Xbv̥*)N����c��嬬k �T���;Ԥ:�bթr3"��UTr/!�!/D~��/��|"Qն�Q��՚�í�V���}��$Ԥ�_�a�w�Xvn6�]wn����Wz�v�H���R���l*_�<
�_�=����{P[��'x;����h6́�k�׉@t_`puR�"����$yQV6p`��82�͖����y�[��hG������)�5��6a�,�	�`���Hggrb/
Iu"W�m�&0w-�h�+|���xa�ˆs��4]�YY}���_���ִ� �	aM�{Bu������m�2L ����爔J8�=ꮪ�c=�"
�(M��Xd� ݌Le�X�u��2Bi��AL�M�m���q9�w@�Z ��86bVߣ|�f�{"r�6PYC�)2�A"o-Ie�����]OX<�:Hnl .A�=�� .��=pa��N�Iޝw��KX$E)�������l��Z4C|���l�NOո����@�U>�	��IJddy�"5n��B���6��^�_!�n��[\.7-�R�;-K@�R��E����R��*Z�T�8���%5��|�]�_�&�ŏ,;��i��4T�����,w�UP�k�/pN1��Kӄ��4� �(�P>�Q����a2�,��Z��-u[�Z�--�L#�ZeЪ�S�2v�;K'��]�������ث���
��C��Q\�¹zĔ�(��@l�֡M��	a��%�G'M�r��I���C�jJ2s�va��������<_��hk�����"�����zw�fkؑ�9�h�y�T2�I �Z�8S�gn�Q�XpW&Y�rn