��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)��<�=�!�7�F�-����8Aʛ��v��	��o�>NO�`��lW�R��)D�w �H��k��C��ݘ ����T�`ڍb�Y����O�GÄB�m��fm������<��޹&)�&���Ԇ��`��^P���
�ԵZ"W*����B!:%�̩s��^x�=�?K/�g�:���,du1�}r#�w�]P�䛗4|H���d�j�_b��0�S�{�^q��+}��j��Â��s��x�5�t�������Թ���(o�<q������"�6Qlc fغ����&e_���6j�t��&�G�(�ay�<�a�s�����pͣJa�e��^���[vd
^��/I�rS��T|P�w������uB���y�j�-J�/����4��L��Jؓ�Y#�<���U1�E29ϔ2���({�-zeRL���օ3+�����`K�H���k$X�E�������P�qO��a�Q]e���+B���1���:8�5�ϙ���� ߸��@�=�MW !:x����=vJ���l�cq+B��&$J�T)�T�=�u;���
ȝ�x��'��k���%r���� �0�'���鲧w4� �.�TA�`@?G�x��96��R3������ռN<��11_aD���v��b�q��9'FNz��΃�Q5����fM���Q�..;*6\}2�� �"U�#�)��e��T$��`�Y_qb�#�vȁ	Џ��E��� 1�0݂��u���%�w���!���ɹ/�Z��Z!����`��
I���zr�(Y��� ��#H�!�g:�I����&ƍ��U�>Ʈ�Aq��4��D^��kF^�|ϯ�|���-�Ԭ����$�,kwc�C���Z%ja�n��5u'2�<o?g�#Ta[��$�*b-{Ɯ��.�P�q����NI�OJ
��+��娡�
��;H.-O.�	B��!��=��T��wع�֨Ӿ�i�J�w��K�i#WU�����h�Z41}3::�N�=���ZQ*	�����]��]y��oK��{�a$��i�t����g�4 +|�솜�����Ķ����˵<�����g�.j��$�Y��KZ�E˻�P�b���&������ND#�^>O�~�j��I�`󕎼Y=2�����GH�i��b�sn��:�JT8U�����Hݵ�s+z�Y��0&�6:�.�%9E��Z�on�p]w8%ݖ�`�������ne�;ZB���ṡ����#xa2�����(��\
��P����)���#$�~�̸����M���<g��<������H�+��m����~�}�<�^��(׏����K�$@ܩ���M����}�h���f�v�GE��sU���I	�>�2�Hay4$������Ȗ���=Dށ�Ś�i�a�[���[p�Ǡ{�
BSn��3K9��i/��WN�f3X��DFi�����,�>�g�@ �l��lZh�#�{ep��1P����DP,wP�W�u�b��2ʜ҂I�
d���yӕo�t|5�_%ss�T�I�F+w+�����p[b6W �!V?��|o�*-�g�ïy�g�~Ԓ�6�����[���>�U��B�S�$f>E!���*8�u3���-)����+v�B��*�Z��ٷ�ƨ�I�B-���n��c\k5i)_��a󨹇QۊQ��V���sR��!,�4��G�����^^�ȃ�a� f�-P�Iy=�+�0c���� ��ĝ�p��&m�.���=����Š�%��Z�0Ǳ�b�x_[�C��nS�,�^x'}O]��E�X(�mdJ:&��	�p��������	�vl�����ɜ���0���ws�;�5ڑ��T���]x���^Z1΋�/�	^��ݐ�χ����7mg`k1�"��R�f.o;��%wE��]O�l��A��i���F�I]� ��m_:��<[�YB.-�`�.o��9E�TZ�%7ʎl��v ��L�| �1	�+�4.��j�P<�d��-{&�b�t9s�gt��h�{)���T�J@�P�4=�]� o���QS�Mw�xy����{��_x:�_R�a��[�@��Q�m�Q�uK�BRa���7�v�e;M&6Z�E�8]�1�P�OA�R����y���U�YDkK\\�NxG���q"FH��ys��g�&Ӊ*�V�3�]\�D���|��Ⱦ�|ރy9�W:��������?/� �fQB��[����.<�C'�ť���C����X'D݀�7\���a�i�T��#m�$�TQ�J�8G�Ϟ��)�LG~wj�$,^�+���\�B���	Yeqw��O�m�pB������&�c�j�0������R37T�m#�5o�J��w�X��<[�A����o�h�L`\yd����2l��R70�uAXj����Άev�66s��g�V���Lb�*I���IF�V`ݔW!�f2=$�a(���}����-:������ �$��k�E�w97̘���>G]�=�`�@*	;O�#�aH���Q�"9�݊���C���?)�$үdϙ`�~t�{���X�����5�����vҢ���x�,�*p?�p�S��z�)A��y�z�x`�~�M����U��vy�������p=w�9[���"2M��ƻB~�ҙ�X�D�����Fm��;X�o��J�m�}����g��W���J+�n�FA@�થ����~�r�4�0��C粃ri? ��%�[K���d���������z��(aI�'��&�V6�7 �1��x��̘��1ٺ�Y��P1���L(���Ы��W�U&r���#Sb���N�,8�l�i��QjJ6�2>|A�G/d�LMз�ǈ�!��L�B2FPAi���U��<�[7.$U�����cQ��86�%�B����K��v,�Nvw�[غN]�	kҐP`-u"���bC���U/'�5[-��E�R��7���Q�B�m���y�ƚ�L��v��lb�z�/�s_��b&����x�RNv�(�ʻ��BJ��/Q2ӧ%��D�@�n�s�Ա�R�tx��,�̈&7F�%�RT����'�-��|&��l](s.I�p�F�qM־���Á$� -ް��6����f����ad����P�ϔ�5ᖄT[�!.�|�-oE�k_�'�ܿ��{/>�7��^�%o��Ϥ1
^FX���u���$W1/a�F��OK}.Әf��-��K���!��V�U+v��pќ��i$�4���u���,�w���/\�����s�)݌o�_�N�ȴ���l]�غY|�f9��ɜ"o�g�����8�Z���hd�YG�b"o�'U5�G��/>�����MWT�mā�*ð���*aYo3ޞ�>;M3�����-�="n"�	�4�
 .��ן����� ���߶'d�u�����Tˠ��E7���DL�L�+
L�@�7�|��������ڬ�
��x����)^a��Mm�yH"�6�;rYH}��Gw�r�jB+��V���ʃ�l�<񡊭զ�Ob��Pv˧pK�J�ʸ,���{2��im��фf�39�#sC�Jm�E��) �9��_���t�8��"f݇Gr�RA{�MoO�ՔSd\�>�
�C�S��N��L� �}���ī.��s��O�`��:��)�����d88(>[e�զADOhb~��_��r�VAb��5ܼ���bl�Vw݁�P���s<�M�-I���U��I	9 +�I{���?�q������ѳvY&/��q�X����k>�y%��D/3f>'/��5f��9�6��wm �S)�z�(�r9M;\W$�/c���Dz2�'��o:TqP`�@��1�+/V��6}v����D�\������Y|��]$S#ɗ�u�Q��s$�i�mm��������Y�e���K��_�7�T��o���gm�l��ĵ��fn���h�K�r"D^W��``��@��>�����@��]A�I�,�����l	v�e+X�;P��/��ǗT�c ����h�f;hOO(�����A���܅ޝ�UB� �$u��u��4[�h���_�"�����1�fL���YK$4���]�����+�����a�#��ntP��;
��}K�*�%؏��9��K. �7%�C�@��׷�*�jfx=D�>����+i�'�]��.�q�;��;�fE	�!�-��r��d]�d�H�`F������ǲ��w���R[�C�2~I��?�|�m��m?�᫢ܼ_s;=�8x��ڰ�%��}���XlI�*�����o9������(��y��m�n�ۗq9�iNu�.fNaoDx�L�]��/iD�U�:���C��BH�CT+`�*S8�MO6�rHKW�æQ�C�s�$, t�_�)6]YXS���,�{R�V7n�`�á߳�00���cZ�+=���)b�qf=� b�y�^�K�H�~ݑ�)a��i
�u"���;���/�JՁm�	���u�)u��n ь͊���������-�ZL(��C��v^�Zm0*W��C�M�x�Ոj�{\�xƋb*z�c�M� l�|�;�F޾��"�d���w�17�R��/�~�?}�)����E���k-O9f$�z1w+��|/3��pV��ے#��#O����y�rǠ�Cx�ң��2�+pXbl��
9�Hh �=���R�L1}�ƃlz�I�r�M:/��0�_��M�5c�Y[�yۅ]P' ���ގIwZ�O+D�=/��,����_��u�\B+NB������2)�ۃ�+?�̜	����:2*�8�ML=k���t�PR%��B�N�Ѐ[TFP@����������U��ᳰ�(q�����E���w4��\�x�$��5�)�F��9�@ȔG�6-���8/�f��5հ[�g99���5\=7�T������aҁA�F�c��{x�0�x�|�_r�=ɀ��ɖ�;��$�!1�����込Bl��p�����.����&��G�LO����;��a�2����x݊�.��>1=�)���yB��
��Kv߭�_quF�P�7���~���o����%Ku��S�:���0}n��
����1�DvZЍ�����c�g�Qm�+,/�N;y,s�s�~�y ��E��Љr{%ɏ�[.gɵ�Kmi3�ؙ��i;��X�4�+2n�	m�h�aN�gb��_C0/$^��=3���U~K��X�>��%G}�?��O��m��O�B�M	z*���k�N�_jh�>ӂL�z��i�V
ڳ�%���R�ߋ�<K�C!�n��=WdS�i�"���	��}��ٚ�(����犤�����	��ً�Mm��iG�a�Let�WEt���=;��6 �1l�M����:����B=b����\����NS��&:�@o�u��gs��?9j�b&(���Y�塂7���D�l�_`�:Q�ձ�&p��7�ڞ2�������"*����1�����r������~�{c�e��Yq� ��[ϳc+^^��i�#���&ș�}ϐ�u�V>,�伃V]��?��[.��7��D"�䂁��{+���F���Z>x9���~��;#��Sq�#䋖ݒ�F�4Bg�\v���Z�9�5�i��YF2.گ"ۤse��q�Y�X�V��(2_üLO��+�Y݅?}�&ko��+�K:?�/��<S��n0�.^���QՐ?���-�h��ZU��B�qe��#Wy��jV5�����!*zE| M�;H�F-6|�҈� S WZ���ޜl!NP��"�^^��"��Adª5RxT/K���ߔ��5!��HM�^i�7?�4>���;=�3��[�b�d�Zt^v��ϼ%Ҁ���􈯾��q�{�>�����O�ܚ�,-5��Ȁ߭��^ڗ�3�%���#�ښ~��$�l��G���u��C����*.�tk�FA�<���nr��.�<�J�>D�޶	����k�	UF�m�j��#��+���Y��<p�b'���d����?E>������e�H��f�>����"�ʇW�V���~��S��R�:���\��?�&�,Yy�|��;V�2�Pc��K7��/���\�sj+3�b�P���au�����.?j_�ʯLr�<r���&#�6�����w!�o�z�+)=�t8E�O3p���E�8�@P��sp���������s2���&���\j������d̓���ړ5�x7�_Ǜr���!��G��6V���@N�LΈ���J�bU�^7�!�d�n����3��W8e���SW��r�M�ګH(��z"��G��`6�9l3+'���B5�;O�r��n����
���6���� E�\��#�jz��4~tܺ(6 Q>�s��2����DYl�=W�$�e5(q�4��VhRa�����7BĊ?P�q����-�&�)�lpI��9������M�!V����]:���<C\�ԱV�Ǥ���5�#c�%v
Z&�C�c����V�V?���6O�}O�R?))�VJ>��,Hԝ�R=fHEh,¤f��'iv�,hif}�7>R(����j� ����������(Dh��'z8z�����a/���S��0�|.X #���"*���ٵF��8�4��"d|�j���i�3�9�3�1¤�D��^@U���zPq?��f�l�o�_�1wEĽ�4�vl�`<����D��R�g��\/Ѹ�p�H{Lz�GZXh��SZLA�XR�[�(�N����S@lt�� r��4	j���$��VU&5�UI�4Zo���ZW�CY��
;�����z�n���]?�DFAS���[�������TĲ�:���q[{�����E΍�r���e\$���U�4bUa��VD'�͌�a�N���ޡ܎��_�]��hW�K�{���8W�Q��	�6�޹-��u�TO�������	���/nd�Z�J��l��4��/�78~����i�c��dc��N��l���;��w;�ƈ?�2 �L�5t�T �z�Ј	N�h�@�Ľ���dyS&��%�kl�]2Q��	���+L�"� Kf6r�v��6TZ�E~� ��z��&�V<�8H��2�`�"Ė}����xWe�ts4S��4dO���8�,���r��V&�`���dEE�&G�C���-A�_����b�Mg'1s�����¦��2�t�`^<��]�#X�" �_�?���(h[A�1��x[�\����Y���S!Y�tE��R�ƶS�4�bn�:d��9�����]M��[P|�& ]��t�Ӂ���N,�흼�����7ʈV_��e&��7V�m�{�l�Q@��a/?1}��-4;��On5�*2G�W�����]��P�%) ���CN��O��k���7xf�Bx��՟	�-���ZѽN3߶���
����\���1@�[�Y^��G�\�S)2�3���D������_P Z�|y�'�9;LUx�Z� ����l��7ԛ���!�M�!ß�<�,6M�0R�0T��]U����,LnӤO��w"��˛m�|��:����W��N0h��.N������r�C�Cu�8���)C��[��'r�ԏ�s5���bl󺿠��(��S���DM��(���@�{�eP��#"Kk�'��P-#��K�����4p��l��|��-/���gk����A�(�*�YF*no���#�e�c,���ɚ��I{\�"|��Q������I�����XK�G���D��/o�橨�'��cXpk�):�%s/2ixY{��!#�Mܵ�=��7^���#Ӽ��g�t}-	 C���Ҵ䜠w�]�U�~ �q��zL�j�Lkm�!C���b����g�t9���G�[%`��?E��l+\�%����0�܀RV1sS����9R-�������D��i��4	>Z�0!D%"D�6�:��GfД�Z���@R���0t��s���4"��O���N�4R�ḅ�,c�;���	�'9 00&
�.�9r�b�G>�~
G�j�F�|�]��r2�毊��ĠH>W9|zc^h�5]@����C0�����-�J$TF,/Z��1mTC�/�A0e�t�±)���#g�is�ϩ�p��P���<��g/I�{��.=g����l,�/HV��:�'���8)Na,'�B���gP�s(��k�ќڈ����~��#߳��Cl���~j.P���5��w�C"�j_K>�Cz��M^��h�"��}�f��>M���k���81�=wd�8�tG�5��7i���|�2D��|\���S{sB�ՠ�+�%��� "hn��1��� J���ӌZF��vn��i��]$NvZ/0��q�%^�v!/}�S��F�.��������J8;x�
9�����a��g"��"��u6*��������uU�^ЮF�D�r���H�.���u_$)��{u��MA�S(5q{�oV����'!�񪅌�� Y���e�+��]X���y3ȁ