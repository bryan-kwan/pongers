��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)��<�=�!�R_酎�����U`�����B��%�y�(���?g��X� 4j����W��K.��xؽ���?M�o�u�m���F����s��f��ȅ�pi6vCUdP���|=�cڴ�3|P
�זnߚ���
?GR�WOpd��I>/A �@L�4�F�]s��1nD��}X:��Dq�m��*3��H����M:�H�b��<�?�5��b"Qn.
����9�9qv��ul;0iWf4�����7�7�5��l����=��0����s��O6���x����L!4-Dύ�O�dJ<�#�N�rN�Hv-�
`���s�Z���M�����Y��'�7��,�����S�J}����k=�<Z�mdT��ܺ�~r0�UoD����%.��0�px�IL��-`.F�xvB�JE��r}��M�*X���}Y]�^��=IRI�T����2�+���˗*QWBG1=a�)��[^D�to��7^��t����D��q���,�1��)�5ߏ.]���V*�aq4O�w�2�
� ���ޟi�JG0���;�z��B���v��c��o��Hg
� Tj�5-e���I�U���@�)�ғ3jH ]0��w��ć0��LK��g����^���'�"9˟�M���f<u&"���%
� *�����쇃j$C�Dc���,[�+Ń=Nz��;�V�Fv��v�}$��d�^O2^�7;�՞m*�q�U����)�	"��Q�Ә�=��3h���D���S����/�u�坕8V��ǥ�A����ְeCϧ�,�V�p*��i���_Ob��_Z��HC���q�s'��9�!�Ҝs��H���ݮn8+{q'[�,-��O���0�{�X"�_8�Ԕ�,�tG퓇̑��Wd>i_��Y�Z�9��k��d*�&��G�W��r�M�_�\C�o��M�*�,��:�%�Q������ԯ�R��K*�ev犻`ݣi���a>}2g��5�x@�q�R^���0��f�DP�F�V2Ә�������"���Qh�5B{V�4�z/�5p�Z�����,�+?y=�X<�=��{�����<k|�o��˔�ѩȚn���@��	}���$���V8��!���XH�D�Y0��z$:aL�-@>�+������a�C�\�B`C�X��!��b��q=f��b���L\�����L٫w�b�&H���'�m�?[��3�cM��Z�E ��Aul�NP���Q��B��}��ޱaNs"��u��N�VSΥ�K�fF�� 9�M]�3	!!GT>�$�0����L��u��7��{)��$6mL��$���dWV�e�cY��[�ԜE��i�=Q'��c�	(�<�t䰹��ɷ2���Av��"LN��nhK�ceP�2F�x������-bK�-��	N	ؐS���fLU����.���P���*t�p��E���n§����4����6)#:�!w�������& �ۃ�>X�(��d�9t�3Y�唺�ML�QB���>�=�-�@>��[�&�0 �~��53]��n΋�@6����
9ӴԻ�Mϖ���`ch��:�@V���VJ��Dj�x{Y�	FZ�V��>�>��4��DX�S�؊��ƛ�#�͛(��%�ڴ�X��q]gHN�#(ө��^��|�Ơ>罓x
J��jc9X���F��oy��rCX<Jj��I�C���֊�x�ݖM��c�/R�lU�W��=A����ގ��MI�k�+Gt�&/�͕+ݳ`,}���C饥3��`{�޶�@q���MЩu<^��"���?�`�7ՠ�@�0�$�Yūm7Ϊt��� h:�2j�n�Hے%�H��jo�=e[+�!j�K�L�*0�ݗø�LV�$����G|��]:�>�Uu����k3�*]cO�g��������m�#�����H:����j�������ŭ��?"3�jN�R���B����&%,�������t�#�e�UK�#/'��,��FI�� �CNK���&�?�-����Őc���~隆Rx��6A8��9|�ur�	���H�c@��t��M�/[�,�������S�48n���+�����$Bx)���JI��ؔC)��)2]o:�܁#V��"݈��6 �k����CRh�q�͜��S<N"9�5��i�hwoO�mn����h���[�:�j�O�Ȗ3P;�G����cO�C��o��%����l>!4�^�h���f�i�0��/��'�Q���##�nG�Ox*���t�Ʉ��kb��;��&d)+J�����0�՞1@�e��o�8&�zv��V�?���D7¼A�{	3	�r�Z�h�̃�@���M�G/�+� :*�Ɵx�Rw���q���|��C�����M�L4;+u%�"b4���9�1Dtox5)M����mtpN��{t{|?�}5��h�/˿�l1�߽� �g���i{M����2��?�e!*~܁P�D�E�N���L_/U�Hh���ߤ�!�{����������!ݔ��G�Ӛ��(��%K��?-ؖ�k��r��SC����8��g�P�A�_���G@/F$�$���W�{�(Jؠ���1�ҧ��
ᇤiq���?��fg"{-S
�0t'z����}A�����7�w�DnFG�����Y���Mы�*��|$�B��^N���jҶ�o	���э�Ѝ��`�4/�?�DS��̧�V�q��KI��z�Bv<�>.�Û8g����"!���\B����PϘ���̉h�K�X9y�T����m`X��,�C��;��D\������1a7ߴ"�t�����&΍�,Zn����Q��?)ܝ�t`̖�k�ho>�=��;b�Ɲ�&����U!v��a��}^����L_���?�ݢ�D<-�_ �� cN�o������B��6a)e�6�F��9^� �����ৱ0�f�2�����s����o�!LyuXֈ+D��T�T0�>&������bUm�L�+:����Ğ<0�ZM�Z�tP��V��o����!�����n�
��!��A�x��Ȟh�V��>���؆�m�<ux-ƞ���C��R%�;�%���B�U�������*~�A�x,����%%��w��%�$z�N��J���uKGm��CA��aQo���D��-��I�	���A�%��YE��TGω�ա��8���7!�\��s���Ð��1��Nj��I��ob�z��T�r��!��]����pv4�|�M'����� �3i��j�GC1�I��{=�`�ߺ&$2��b��D�')
/G7C��?b��B���Is�n2$�ؑ		ц��y�#��0�c�K��\���q[�Đ�m�м�����?a+?͘Ǿܕ�mЯD38�⾕�s�9%��F�J�����6���M���6�qPEҟ�����!��|}~�߁��m�;������\��X�Sm���t���0R���|9~Ǔۻ]n��u��Y���.g ��K>���m��u⭰I�V �4D'-Ǩ�Wߢ�����N���7�7Q�����.��Z1̶&K�-Vԩ����rX݉?+q�\�*J�3��z׋�J�	���dѡ�+������k�x�Z�8���Q�]?�.�>"`��Dm�s=h�d�6fN��j"�"dLH*�-��p�T)t?�],	�A��b�b������<: om�;��֧Qc�-.��m�t�O8�\��b�SqNT�;������$��)��9�*�7�	��b+R�*a�0cG���%�U���f�,>�<�`h�������Ʈ��|nv�����+�f�%����:��6���LrT�lS��Ng�up�h������r� /�W�_<a��J� ࿡o��S�#?�i,2�D�$5����cN1���S�r��t-zSd��tț�'�*]�R��.�oB�,9^u��q���4��]�#5��P�齝8��D�&j��%M�tw���NM�r�>䫴�U�3��ک�M%p��k�lC�i����\!Ռ,ҽ��u��D���D�<�C>�	�ꐪ�Z=1��H��*��=t ?F�����Az��_���p��0�9����rK<�[�	'�⼘�X����Gnf�鬆��\>ae[Km`-�J�E!kl�Ddf+�VH@,h��P������p�'6�V*�|k�H����;�Ź�������㙫�Đ��y-L=�ũ7�����5�=M'�
O��,����`*OWN�$L�4+L8ɹ��@%_��20������E���U8"�>;Փ4���q&e�q���4�\$�^����y�Sa�pv������������U�_�$�"{ϖ+؎Z.�g��L��zU��h�~YeB��-(+M�=gv�o�'��%��d�
zi�vĊ )�����A�˶�ꈶ,�7�s��rF[��4���8��H���&­
J�Ç��l���عlђ%���4��2���r�x�7<�G�3j�!� Z�0�r��	�cZ���49�?�P��R��[{Fy����"�í�4>����N��|�94q���;�
+R��ԏY�\f�B��+�����h�߬�*֭�&L&�0�y��[�Ց��{�MˁK/��N�d�0Q`��#���*w�%��H�z���Υ/��50c��Z�MM��K2{z���^�*�>� �?�K�BN�_3Eh<~i�c�28� iJ;�6�r��HP_Ϛ&¤���Y$Sck����D�Mb�n���u�)�5�O�m�6�F�:L��<���9*3���!`��d���F�q�sв�|��ۗ�{�̘;d�n�����-Y��;&u�d���꟟FS��ܠ��
c�T�Oe�g|f�~v�W1�Ǿ@��1W��)��0P���@AYeSܳ	�{�b�'���/6�S�蝔=Y��$�w<��vfX�H�@�lV�e}��� ��1:���q�Ҩ�W?��X6ր_j�A�9ʛ�̣�q�%���Ee��=&*��������?]�~΀k����*�|(�U[�y�ΜJJ/L"��T�A��ϮJ;Sa1�4>0�RG�ɐW�I� �*�L(��Z��#���VHC��42S%	C�-d���p��9��
u��>�t���ĺ��'��_�?���^�1V��BB4*I�X��W�2�M��Zk���בn��\��yw�J��֋Z�*B�5��j�������0R�34Ԏx��Y��h��@�t8%�?2�b1�f	,�=�"ҏfZ�WR@kw�8��kUCg���j��w^|.s7	]�ſc��&4ο_,�T�g���
���Q��*�Y��L����q�Sus�� A�$���bSY)o���ｨ}��R�l�Qۖ��s������v�z:�t�@J�hX3Р��Wo8�P"�h�5�PD-ӿQ��Ic7X����&B������f(�������b:�DI�V�Ֆ����m^W!��\i�lEYU�\��2tN�H�
cʁ�38ɷi�Ҳ��M�5�oQîjO7M.�q�d$�;:3E6KO��<r�G���8N�	+SU`FYt�v �4mS�Kt�w�R���;j��c���.jfY|���N���ς��-���N�%a��S1��ŏ%�YH��Ux��[϶�|����+>q�?T��W���m/���$�J$ ��CZ����CU���k�KG�eEۨ�9/W�B���H�$�9�k�������,��'<뉵�KE�r�����n�A!�S�EA�B��2Z�\p�T��ɬ�3:r�����[x����=4�����:�0nN��6{������:�@�M�;�����r��N�FD�i�9	�gt�⹾++�=��7�Z�[��=~b�����(|�XA6
��_���CƈI<��묷��M��>�<����8��B��yO.�cO>��E�z��Z���<X����z�8J��NkM� d��c������/���=`�$rJ�s� �����ˢz��3�U�>�u�FGQz1��B�`_YI��A���� K�c$����]���Y�@�f��]a"Qy?�� �>��aJcqyv�}{a�����݀�!DϏ.��#������w#��@�5�O�roz���NR��	=a2�B" �`�o1+-�O����G)E����5�L7d�N��K^�c�4b��܉ǏJM�1��ԚC�'�+[�� ���>��~�g��!e�.�Aw\A��5
mQ��0C����"���ސ�g�H WZ��#�r^ꃡP����}��/j$�I��!�-�����1�|琉#�|��|��~7��H�;䀼�8��"g�֨<��Kg�7EE��,%kz�����A]����}}g�k��z���O�6E� ۳3o�;V���+��)�ZT���a�2�t7���U�������s�/XU� [����O�����=��d���1잠���ym���w�4b|���m����/	F����Q��U�HO!�	w<�����|N<�SQ�U��_�x�wr���C&��u�����صܨ� �a2E)O��Fv��u�(�v�^$��[��ٻa	�������*|{�5�._&ă�_��	<HqvN��[*[1�0��g�r�m�x[&����p�7�.�4{L�W�K���z�T0��+�|zF]`��E��n{��}|�:��~79���"��6�z6�	�(��Ux�n�ӂ�0P	o��r��0���O�BW��l�9��(IV3�Y��vM԰^٦�Ǥr��d�~<���~x�LSEq>�Afm��q#���j�ʊ���]j�'s=�:���ߘ��ܵe`�.3��~h?]��ַ����+�b�,;Ƕ5)�Q��h�b�-�)*�d-a�N���̻���1^���@���Yb��ۘgmR|�b�-��Q$�st��G�]-<$+�����{��r��f�r򑸰0�&$H��/q��$��O.���O؃~A�H.3���ya0^(s������ߓ f����k`6���g�U�� �N��V�г^��
�eʳ��wR�:lz9p��)*�����#S7�i������,�ڗo�∬��(���R��7����`Ch�g��t�Z�cX�c�I[H����_ &Z���*YH]�"�~�܅�s�c�7Yu��D f�l%������#e�~�KC�ުN_�ZFt�4��ʎخ��z�y�2ޢ�ʑ�x�a�v
,���w��}u����SgQi�G�T���'�J/�t)���G��4]Q*���X��U�����b�
�ָF*Y�P��\�d�wi��+�M�k��6�65v
�&d���,B�ȼ�p��˟�2
6�\������R���a��z�l�kX�!�f���<\z�w��
E�u{�d��@�*!��qͅK���T�����<;=O�ΐaPЅ�O��@;�©���>4-���Ig���7��Cu��p'y��zgC�A���a�F�<��N��t���"�S���?w�wx�V%���:� ��I~F��ᣋ��i���N�W����=�j�$O�l��A�̕��ŜqG1D��9�Oh�]�r��ߒ�i�2RF�w@����Oݟj;7���'��rB�Q�z.R�&�n��8�iɔ�\i�T�`K�
�o���_����^P�;�&<#���N�-[ ��PЉBa�)5�\���uP晜v�ݴe��Ֆ,��!1�;:��l�=9�Xc�W�[(;�y<O����oS�Õ��>��
�S�V�@�W#l��h� ���K�<��ǂ��nQ}ml�������NcK�I
8Y1i�@i�Eَh��k�QO���ͺl	�l+M���l��t/�(����'��
Y����Gml ��:E�K��ٿ^��["��p���\P{��{r2}����ba1����MhdKb�S��O�xf��-��l����Y�Z����.3�[_k��+�cXa#lkt���z�cC1��N	v���Bќ�B4���.�q���<	��e��Y#����1��U,h��h�0n�AߡxVH�'h>Z燬��U�-�a��w�1Y����̴Ts� ;�?:�7�B��͉��I��À�ysn�s��g�:�����Ǳ�Qvsyxt׾�	�+A+���?�ǧ�3��ߦ�K�	�nk������h�0_�W�׫�U��]D�e�l%A8�H��10�4#���.�;���\)��A������n\=|�6� �D�e�X�����o%?SCG�M�3°<�0c�_��3��N�-(^A:�W���r��و�v�.ǼkкEe+��o�������c@��ڝ選�d�x着�b^b�x������Hfbu.��Av�(�j��iԽ�{��@}��g��L6�6a&R�7V� ���~^��� ��Vd˸>u�i8�p�₟I� |:���W��	,����p�&;��9�h;��M�vU��
(��T�Ds�W�?��g}�^y<q�����K��i�D ���&��G��u2?d�����rK�= ��s��[tn�����G�d8�j~n���� )�x(��h�\d�S�Y���<'��q���X�ns#s���?��I������-��~�a.lǳg�(�ƴ����]��nnu&���� ���?ls�����J�Ѯހ���v������#���)�I��4��})��-��D�[H�x-E���S�'�B���Ǹɵb�L�N� X�`H�W� ���DM�j\����aZ �*�l�A!q�n�1`�Dn��i�N��9�!S�'ˏO�8L�i��6�l�`�U܇Ԣ�����'*x(������oo=G�3׊��*�7���-<�rv;�S������	������d��á�t)�����"?%�Gnǘ�a5������ʡ�n� �![ �z	��'���3q��a�޴�ŋ����[Mb�
�&��5�*r'l �؞2^��g1�(��,�Hɪ^�O^b�Z�k��_f)\�k�)��q���Z���d�"��b�����_{�^U��ک�䅊���
J#ٲP%\�*��a���"z��d�*�x�0O��}��)Z\�}<W�p���S%qf�cQ%��'�m��39+x"��?FX�%Lz�%�J�
�?�y@�����E�#3��؜�v&y���N����RA��S�9��-���{����v�U"Ѐ�=�0��6�@��^Sᡑ��Ly�L/@�b���,c'"�`�{9n^�cc���k�I[�Z�F�,�$!G�@M2�Opr���:۱$Ո>�MQ׫7���
,�g�0�M�d��~�b@&=	�v�U�ì�����A݋��/�7e��W3p��ڛ�6�A�N�_iL�^O��I_QX�6�� T랐��Y�?ˮs}�e���q��<h�Q�����@MK$(�%�C�ɤ�2�����A��ܽ�m[v�m�݋y����Cª3����'Y�ҎC�o�A�c�]��k�P0��v��֋#*����V���L� �&|��<o��\������H�� q��`��g��#����=El�؁��BM`P'��16a)��+/��{���_�r��>���AoX0���(���59ݮ���S<x�ZS�����m�]�8�l)d�Tt��5����?Kzc�%'��l-�k{60�O�z�H�ӵQ� [�s�.��?��n��ʫ?�?#M�.����;��qq�6 ��!��o��'�`IH!+�lL;J�hbŊ�DV-C�C��NP2J�TJ88Dߗ�6�� �T�D��ߩh���h��=Z���SK�SR
%��p�ߖT��h� �y�ɤBR��V���%3�Bhn��}w;\��~���BP��8����g�`���[��~�l酤S�K|(��9��/�D8I��2�N����f��>csY�Ax�T�C"��P3�X��ܞ�À4��DoQ�e�*i�1�6;�ٜ�F�#�
��,�+��c~K��z�޵-�86�T�Y���n�ɝ�0�.x����{�YQ����� 
�4�/s	n6�nNT5D�k>3������W
G@~V����V����\��2\�*WA4�fiB�
��q��`�*O�JeB����Ҁ,1����/^�Ӊ�q��gU�da�Y����38{hg� ��ȼ<�]��룐�M���3�2��'���g�B�M��g f�:�<	oј��# '�>ժ�Y�!��r�Ҍ���#�iD~��fik!��N32-Hl����(@4�\��0M�7D�U�w�*<f�ݚ{+�^��S�V)�[����*�׾N% �5����FDٞ�I���~Ϛ2-�·k�e������s2_��~�j|�8�׶���� ���륡Z9-`��������x��(��-���O��"�꓋���#aA(7�d�!󡂕�d^H/� 7'w�0	�d& oS�]u�����?�D�فDEX��w� �DBN�H�;.��A;��x�6!�9xt�y���Vo�^
'�7�q' �nE�-e0�����=m�|��7�vy0������c�=`�د4o��!�wm��9D�]]��I+;5���T/EqE�t�r����2�}u�"��b߲M"m>��b�lDS�;��}���W m���b�6�5��na^k�����i/ͤ���bVY��u��v�O��I(��Kb��P��Y[��(�P��e�����l�4i�i:Gj�
���|W$�{5�s�3Et{���6ab�
!4� �@)]\���;啲2o/��m�}x�4P�jڙ%Є��F߇��>#���t���/!�1��|\��yf��e�j��0��x�i�b�NF+hI����.��ꏜ���u`7Y]�\r�g�vG5����ɪ��i��2Z$�$��N�Mx�>��B�(�w�li}�\(zWn�H�'=��%�Lr��&���W�-_ɐi�� ���	:�{���s�
O��������fs��M�	��� ���)�:�YA��8?N���������� 2o.�O�>Q�f9������
\~{%�Nr	$�'�Y&a.�4�°�"���_#6�l7�^��%�yItm�EQ)��Ɉ���ONK��2 ɕ��-�ɥ�<��g���ɤ7jf�I#:\���yiOm����F�J]?��&�ti�	J>��C�q�J? sP��[�l������_��u`X�R6[�p���:9�sx7�����	����8̲���R��~��Q�4k��&��_�za��-A��#I@�Қ����q��6r�ɓ��-�ϡ={�gH���y��c�g��������lʬ��#0�u�<Ԅ�l^4�=,�C��8�#3P�Rp%ƶ�~G�8�ٗ#P���_w��,H���ci�U���X]��/��R�M�y�nפF�
�CNQ�g ���'b�ǲ��X0�:PχD�r�r��y��틹�P�G_�t8p��T�����"�˛��)��u�z��ߗ�?G�x�Zo�79sR����V�����D�S@6�p��T�%#���ep[k��d#�oS��y냷�6-�9� z�/_�s�7�Ev��D�l�R7]o��L�)v�2�WI�&��Bk�To�N�a�~:���ӫ��Np�u��'�SV��{��|O���A��4�j�We��Q�O�J�0A�؅A0F�?ۤ\��M.B�A!r1<��Ao4�V�-�]Kȳ~Ф�%�>~�	��'$�s�p��6�s�W��r�o9i8�@�=����R�ʴP�h<0(�h\��$����T�fA���Xt�Y�;#f�C�x��B��<�Ca�&zbڃhZ@z��Br���"U?$�+~�n�I��|n=�:/�B�j�LSH��^�#;ʨ�%1�Y�Tvk��t��n�Μ�^���ו�U+!<��o�Y�ne6q��k��L�ӗ,���*&�Mk/�5�C(�o@ح�hNJ�XPv�X�tm�٩D+��fO��fV1����'���s��=[�.v��E)��d�S=�Ъh��[b��Xb�i���]X��Uϣ�'�+�"�-"�lL����UE3���% _��������]���2:���d��'#:?`�������V���|c䣘rJ�|\bAaO���GPE���q"ʩ[������UΝ����&��0˪g�A�����R�hF���~ �P'���2C���;cKIۍ�yЇs{c&(L�3�]y���1�	�{)^\�ނ)�b��UA�����6ye��rٕ�� ;��� ���8�LCS���uLH��v��|%n-0vI�i2�����`[��U��Oe�˞�/K��X]v>Io��&=7�8��*��Nu��T
n�ح��)���Vl�f�W'�������۟M�`Q ���.l^����������I{1JڀQ�Lm�d扉'�km���izһ�Ӣ7�KLD��w������em�(�ﲁ�9�[�d^��>�`z��
��'��o�S��vd�ݰ��*����+h�rZȲ�O$͏�!1�9Y@�J��d�O�M�M��h(yc��C�K��*@m���e��(E���7\��)�)�;��-��Y9��8��0�.�����?���ރ��y�3�ևك�Ԥs2|e��¶�G���HH[&����Y>�'E]I+�d�l^���43����Ŀ�1�b�n��G4�gs�,O�����˦O��O�-Y%���k�>m��צON���]��`����p���2_�2%W_�JJ�;}E(���V�����"6�B��j�c�6X���?t Zf��]	T���!]`�����R-���aX�q<;E���jkqZSu�����[hk�(�G�dv�Ϝ�pa�sT���ć��%���Ƈ�.s-�Y��2����\�1�ah�]�]�%���8o�+!oӚH��5o��Mޤ��Jf�i�!�b�Z�؇Fq�C���#.=�έs�;�4��ZKO�$�D�F�#���f5-�-�&�2^��ab���p@�-�,?4�?|1t�L{c��Mf-�w��M��0�vM:��iՒU�,�=?$H�ՄL=9@K�M�Y`U�pn�j֊��_eٷ�6��x���7����{O#:Ð��X�̭�~��!@g/��w��z�dM�w�<�L����&���z������_�1k�4�|d#��P&MF��g���w"?�l0׍�IͶ2���F>+�mM�2�IoA�[��S@�U~�$��C���DGvƋ��[;b�SN4A��/���].�1��Y�|ho�nƉh����&�(G��N3�V��դK3-���u�����EBz�O���pN�����(YٚzTD�~��%,Q��~bc�p���Q�#�<��=��jF�u��������oK�:�/�/&�>쓉�$�U�GGf��6��Bష���7H��J%������/��iؗ�py��Ę��.Y}LS! I�p!��ُ��Bd@	
ж,(\�=�W=9�'od�L�Hm�M�<��4�͕��B&,���N�t#�f6b�B�]RY9>P��1�<%s8"+��q��z͗�A0*\�v 18u��O��!F۸M�g��dgǷ�T�?��e���pN�A�m�I"$��5�3<(R���e�aV^���`���",�N#��26���w�<:���a}t�D�1s��3���*S��֓n"���!�k(����)+>ȋĮ
��q?eڞ�V�@@R��#���HS\�6����fls�2F�:��/T��!3����zHX��o��=�{�L�e��5PNs�����"�(g�C<h�(y�b�!u%���UD(����/������*nØ��(NGu|�Y�f�>4��V��q4���U^��W�LP�Lz��Mr�pSs�'�1ͼ����h�&ޅ�����ڭ��`HXrԷ*h���#�}�;�( D�D��'>�|�H�ӟl���EDP����B����-#�f��'Cюu��;��[ŉ����W7{�B��.dȉ����^��ᗝ}gr�!�cӕ�V=K�UK�R'֚��yg�}ׄ�v/�����'A�N�	�Çhӷ�,6.�
 _i��Rb���&���$16K��_͓��Ą*�(��J%�0{�z�y�z�����+��c
7}7��e�}AC�ƌ6�mx���!	j����>�y7ale�x��8�޽Z�v-�FǼ�QV�������m��uc����`^����o���_���Ă4�ǺrH�aCc2\Gx�_���5,��L��'��C%i=�`�V7�J�%�KE�2�kq-�Z��wC钬��G��b�rr���mp6���ƽ��
 �Fb�.`v*��9�e��E����3Z�?X�*�(�{��~o,Տ�#�\ ;�}/�ʤl��>��"<s�����%p��8��(#��+��ʭʊ�	Z�r���;�%T��
e�?�U�[�a�Y�@=~�կ���'B�M2��ņ��i�p6��b1�~'5k�Vۯ/��a��I#�hE�a ��j5繑A��XA��1C/[h�K���Ys-I�_�o�⇠{��B�Jl*|�`��p�0t&e	�2g�(m��K
�;��*�ӽ��3��YvPnIC�r��zq�O/zlQ��+j�=��7��;GW� ��&�S
6����b���ud�4�����N�!M�De�C8s�r
���c��Z Ke�#V}ʮW4^�!4c]���|2Ѳ�X�"�����h,_J�����.W_�ו6�%����A�P꨻);�0x��mc_[v਒��&�ayl�Ru`�M-�a<1�G���L���=rP�d�=R0�������V�z��Ǩ�>؆��S�^�	����^i����j�ϛ��X��E& �@gנL����WDf,�Uemi�9?�qaz���o��[V�ᛣ%�z�a���%�45!� �	�j��~/A�	�0=S�~���
2ߺ���ޯ���7r�p�zPm�YU��*<����>.Q�X��p\�!�����e�J��$�س��6~7�S���ԞmT�+�?*]�����M�b���5��t�Mu�{̂���Ў� �i_J��C����=J��'��%�W��2`��/�tf�t���`ϊ���Q��R�4
H��%�g=�DK�|��n�X�="��|>@�	͎e{F$Z]�%j����*�e�)���>�=z�����֬�N�:?}