module song
 (input logic clk,
				  reset_n,
  output logic [11:0] milisec,
  output logic [9:0]	note);
					
always_comb begin

note = 10'b0000000000;
milisec = 500;


		
	
		
		
end

endmodule