��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)��<�=�!��PE���-d�M�/t�v��<���[h�dZ��M�O��#���UH����;�<��`�_x_,Y߷�u��$�ݥ3^�|��Ō/�E�3�|To���'�{^Cެ��[��ǂ��+l�;�{��ԏ��
�d��,?����V���D:����@b�Np��
-� ���An*|����?&��"g5T���tl�h��Ն��Gr�5�T^c��`��TО��&^�fQ�k�!kw��̕��v�-":�7
H�D]���C�F���	���R2�����Z̓�J3ߥ�� BN*��_8����K�\�c��Z~It�sC����XQB�m[�����Eti�:.n���� ^J*.K��i��~P1�~����H�a�"�[������/�F�j�dw1HT�̰X�x	�4��t!��`��֬WA�dd�x��0��f �)S^OY��"�	j"=5��R�ԦU���b��=�Ix"�i�TP>�W�@,鵒�3r	m$�� 鳽��qó��vr�AaVk��_T�9Gz�\�M�9$��Ω$�w���;�{�6O�H��Ud��Q:6����6rY%
�.P���z�g� ��J挷N���O���"�����=��/G�.j�Peb��A\�{>< �q�X�^� C���_"�}%�Ϸ�����<1�@X�@A9\���3Io3&�´�<�>G?ڰ�+件��ye����k���0�F�5�qtyI��@K �u���|��:�7�':A�m�.�N��g=��`���;��7�_=N�~���eOZ�� "P���tHۯU�F����%����Ěɞ{��;n�ig7�}�3[�.�����j��|� �e��Y�C����n��n!�R���&O7=-D0Q�i���Q#�ǤS����s�84�i��R6��"t
��H�b��aNwnE�"��e�ܕ���OGR���,��5u_TNXG�M�>;KYb��0D�{
i�MWYa	�~�,G�߉�qd ��3����� ߜ	�s��{@�[���GJF�;ܧ[,�k���}87�T�h9{���#T��1F����tp)���5�����EŔ+����_���� �T��Q����t��G�K�BgZ��Zut-��],G���c�k���G�
�|?K����Ȃ�ncE�8�5(�"����u���}n��W��&LЖ�gL�{�`�8g���\� �.�� �/��.�?�]\���2��I�t�9�Jn�h�84�yk\�H1������N��+	VDea3���!���Ҥ�����`L��E�^���|��/�"v�a|�����.1�r.D�Kt,�~��dŹ^v�w3װ|�5j�����Ս�8�v����;b<B3����p ��A��ˣ8��F��+!�ڣA]/�R3�����gz����z������ψ[J�@�/E\����y�K�}M/p������`b$'<�V��)jf�r�.)���#�����nha���LuB{n��Fӭl�K�X�KHgh��a%�9�6�{���(_2�5�b?2 ��N��~c�o<�ED�o�ld\��$4k��S�}j6�B��=���4�f����wh���[c
��.<�Ȱln'�����0�Ѯ���@ԝb�+u���\�w�����7��S�A1�o��~ȝ/)�/X���)@��O;�v��F���\�^O�!߀h���2��)ݿ47: �f�Ɲ�}E��>��+��i;j��;�m��k��Ղ�=�x���׻�k�с�F�vM������?��û�����7�zE�Ң�2
G�_�������xl�V�U�Dj�;���٢GF#�1�aI���
A������M+dD�0�z\ZV�	@�2��u�@~g�ٛX��>%�����C:��z��wh�6���i��&�&�p����黬|	����0�X=��v��W�f�v3��<��X�$�.�g���|�u�=.����� ΤXV�W��ɲ`.�`oI��p�^#�5)��4JǍ��g3����d�6�$aT#>�!������eUm�xy%[GE���e�5�x��_�� �I�̭�Y�=%"�L[ҩD�#�Q;|�nB�tA��h"5�?8�ߧ�V=��7�^��c����͘���`ť8vP���M�`�'S~|�%^�͈���(ʄ;zb�	QJ �s-�Kw.E���0