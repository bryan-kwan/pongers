��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)�2������2p|�t����9)|����M����~��/���z�����h��ut�K�5;�5ɂ��٘��Xc��~�x�?N~{�)���ˮD�0{cV�d�m�8�Z��ͩ�1��|��if���9k��SH�Ɉ:\]>�6Rn���p��E,�	UQ�� �ʼO�a�T�NXÞt���e�b�"�M������uB� ��d)�q#�2%���d�7��1���$��[�e���忢���lW�y^ʭ��S���U�<i���5��`�fkc��S�}�8G=������Ѵy�"�'�]i�ݑ L��N��o�{*���,C�)�Y�KN��~u�]��D�����T���+�G/i�%p�A�ώ�ա����{sB��=���͆�ِ�ƿ��-R�$S��dKG�����4�"ma�j��	��rQ�(��a��V1���}\0��P�$��H���SG�%;n2%Vv����ұ#Gb��1F��ٺ�;�t�w��A`A��T���o����8���l¡w0�~�����Q�-F���߼7��$^���[������ȼ	-��	<�)Z���tM��=<k������"��¸���Uӫ.���~�0��f9.�e��&��o�����U��.��G0H�;�O2x$aZ�BkS��Œ�_w[J�cq&ބI�� n*��{4��vs��Ob�=��s�~�>��U+,%��}t@�|Wu<x�GFe*�a�t_`D��ctJ@ѓ�T7`-�;Ө��=8���RI���gM{�>�ս[�2�ľ�̰�g�����'��g���m�����;n��4Y�K���I�w	�)y���x4�Q��p���u�ݮ|{��L߽�����^��Q4�,L��`������� 6��=��Ż��P:Ƃ���)c���c��򸞓^5����-$�D��6�V	{���~	�z:$l���WS$�a!��qʤ�Ź�>��u
7:��J0<<��E� Jv�W�-h�^������zS�|	���0!3O�@^!.�K�c|�,�vL�+�S=�C�L�-!-Y|�8	�i�=�Y���y6�\�V���R/N	6�\.,���2��̮��y 6��{���pW}Fz�[Iz�=��:-Ϲ����2|�]u���<��+�������#����TH����������x[S�DGit�sgc$TCP?�Ւ���e���k�� �[;�E��iI����m��h��1-��k�*w���E�����
Y	�쓍���I,�-^�ԧ7�J�M>�+p�׫HR����;U9s�����jVh�s�9=.<BB�LC;�����U:r>����1l�[�oX���i��ү&��X媊�8j��è��R��M1�9��Q���^�VL�[N���+*ಹ�|�#���|���!>�ul��)�7amxi��#����C�GX�Zi��1�J^��3ހ�䎟����k��
��,��S������?@�`���2�U�t��YĐ�:�S� 1L!��%���F��Z2�	������jb�F����Nv(}o����x��C�f:��:Έ˸�g��41�5�&��7��tΕq_��a�������F��z\sҮt�eEFeR�47��tO��aU�� Ն�^���S;���{��W݌H�B�җ��,ܻ�����=����p��bRB˰'�_ƽ�\Um��y ���G\v�_l_˟z���%�{�=�U]&k��ƻ���A)���ٌ9�B�Z�}"q�Z1����y��δV�b�!�� a6�a���I�ø����Ԫt#�zV9 ���D/^�W}?G
���`�@�.}Lr���'Q�_�$5N�)X\��V���$��3$��{���8B�9��?n�Q�Jn����A'�q�o�s:�e�q�/��6�����$�����x�.QJ+�ku>J�Z��&ÙOTJb��1�c�<�n�Y���5w������w���Lm׻�؂�A�:.��A�hS����9���KŠ�g=�h��0L�𛝯�)����������c�V�?�qj3�֜����eN�$�J�/�X��YY#wuR��n>�t��{���|IF E����Dc �"��xk�K_B[j��XF@l˛��O�7��Z�P�kF��G�߹�`��g�0����֘A.���6Dc�	�GW�޸X3P�@��]0'4
ȹͅ���;]�õ���Pq��Ľ�-��k��5�L�	�A�sw`'���RSE���-�t���BSb��2Qn���&R���b'��`����`���8�6�O��Qh�������$2Rz�`r��p�-��	�O�[��8�m�����_�7�Դ��wu8��������������w�R��y�Ë&p�O�P���/d�S!X�t����~��~W�e�k��;�oS���wm�8���ȶ��paaL`KȨ�cNd^|e:moj�{�<E o���A�F�����s� 2�L=FUPoYР4��eP:𪂇{:� �>:f�`����jM�:l�V	�W;��:'_>�)�y]�� ]�<[ ��AY�|�Ԁ�v?S�7"��
�<�ͧ#��낚�P��{��Ϝ��߅n�i�l��D� ��>p�ŏ�\�)�ָ��_f���đǞ���q]�~��QЁF�kj�`8tqr}w;�`��c�4�C�r�O��'�	K\�2��u<�X�A���5l`�G�k�L��Cw��B�����F�`�t��^Ii�:�^�
ہ��ñ�v�rS�?ќ��YrKU���"� &�m��Ս=�!�(�G�T�X�8Oc��_ ׆5�:���0P�������6g�vQs��=�/R0y��bg���jǿ|�❍�^p��=��x�)�=�$���=�j��@�y�z@m�-��v �x�ţ��6�߅_����%�"/�w�}�qА�3�'p�����i��~�h:J��E�t��֛��-�u՛�,!���f�%��qg�;�8����u�DN�o\ڍ����@�6��k�UP�Rzq�3�د�"+�b��j���)�16
[s=M��J͒�J�Mi�"�-]�"��cd6�G��'5���H�l�a>8�'���#c	�ra���Ֆ��-�%�Mݵ0&���9t����x?�N�W ut���WB�IU�����!bs&)���w��}n�f?޿s�6��Jԡ�*j~��*�n�K���� �+�T�w�Hb�w�C�����݆��U�!5I9���*8�e?f�`6�$;��^�T�+��)����'U,�z�Ŵk�`ͤ��	�ALaܙ,�����L6�F��}�k�B�=?EW��`[�,����u����ؗ^�i�t3������<��a���*;���!��-:�=�l��,�e��i�g�ػt��6�~�����>��Ċ�A�@��ߴ�̦�@>��Ѥ���K�~��7x��zHf�ʠ��
��9��~�@e��H���"."����Õ�Z�g���c���nqwyA�V��+�°��t�9��+c,yH�m.�	s&����d�qG���\{�g�P�!��D����)�����c�Ɖ�93@[�V���5�b'��/8�|��(��T���\�,#v�X��g�� ����x�V���ν��r&+��~�z������B���."�Q6Ä�E52�?+V��g��[�%q���i�}���'�l��inS����F����-"�tk�m��isY{o����x����ؤ�:�?�m�a� ��{)��Lԋ,�X֧C�q�`A느���`2Rt�'NVB�%���- (�LŊ��N�>l��O�^��L ��r9��q�]I:�5��n��TW?F�7ٛ�P֛pN���/��%L�K׬e߿�E�by*9n�!����X:��3k�:闤>�-?v�[4���(8��x8�d��A��v�*#Pj]���=�4!6?S����m.C^O�����o�v��l�W�a�N�,���9�4T�*���h�	��a�]��6���:������
����{wt�-�h�9�y�'%�5����N�U~�h_�T�q�j,(��>���DA�U&4�Pq!�=q�ud�����ͦ��P���R�J�l�
�����~g�5T��N�V�l/\|���`Fa`�Q�#&x���uS�oߛlW�3�Q}�����C�����R.Rz-s���2~\V��(V3C�@�Qc�!-�;P��, �l��
N���پ�k���ݔF��'p#�\W:�}F�z-X!dk.��`�Q����߇�>_��/*���Tp
�$���ڇç�0�aBD�\���O>B�.؄���Z5��2����2��p���T��$5RW�tfؤ��x_����;m6.H4*�nGIׯ�~3���ֽ�D0����p�hʬ��D�,G#2�mdЧH�7�0XM�t�H�[<5�,%��gύe%"��ﯮ�������ZA]���h?{.=Ɓ*]�5
��Kt��r��L�5�� 6>r�QgW-,�!�15�	�_�Y� N�4���IbF�Ӫ:����;�]%��-:]d?� �8J�'b����b+�+sŖib,kx�DW6yƯ�D����h���!���a~�`m�X�����k�܈v�y����'�-<�� ���$�,Ԝ��ʛ����`'zz|߄��2��K�L̹�>���9#/I'��u�UcTm7�|!3z2(�7n�x6���vaK��ej��E����C�v�Fa]c��g�
w�؎5m�)�1 ��G�����KXP�i׹8RWn(us�����IGf3 �Ɩ=!��p��t_1欹�=c������V��J��xs����:���"=9��`@&��>i.�y}v��O�����v�o�8U:.Nq�K��a���$#�H�����\�֎Ҕ</1��s�͖[���zy)dY��O(*�F���g ���uʿ!�fd�O�F���<b��+x�i���da�YoJS�N��q�_���-��Y�B������s��k {��E綬��N�5 o��,Z��:��A�K ڎ[$��>x��6��ҥ)����qo������_3�Vߌ@\�DoD���^ѩ#��R��t�l�����
	^.�٥N�v���$�!a��(vp��-�\z� C(]e{�2�O��b��F1h�1�(A�T�kwk%^���Q˔����Wf>Ȅ�cT{ѝ��YX���+�r49=jM yՏ�mF���Z.Y;��>���`���R�c=��E�{p�(k��v�݅�+��C��)�"�K4��q�`="L��W�=�B���jD�j{�9���<�����p3�h�o�vL�Q�^�[���ޠ�F�G���U啀P����$��zkN(��(HiUJ�I��X�P�PS2l����s����v2�ȃwn��a9˯@8#��w�H�,J՛m۝��Q��	�$�L�k��G	6�	�nT���ڭ�(�P1�52��1㮿�FS�gB��$�y%�(|����M�J eU�,�h*�Z�e��Z�aM��<j�1�O�F-R.�}]�F"����#EvLpb�dԗ��}]ċ:rհ�C緱���g�)��h�AV	�)�����1P��Y���ὣ���D�ӏe� ���k�������L�^�p��ɶ�D�Ȯ����A>�T�j�i�%7A���+��ֈ|�1��8�RKEe�a�=�J�i���=�Y��M�U����b���s���	���~?�3�1����cp�B����Eno,%d:r�,��-�]9�hh�>��3��Y�4��+�Eގ��8��;���Ϋ���q�jQH�(r��q�J�X�.�Qۃ�e�նetE���w�E�_K���GWJ���v�4/��ⷲ����B`�"߭��*e��cƳ$�k�읳M4׬�߯��P#@�K6�;D� ��"H+�[s�1�/I���af��.= N^BM̕_����*����Y�!�|X���C�^z�J��i��>'R�������.�аe|�3Y���
�`GCN�	f�H� �If=��pْqb��Ęu��%��VH~��^^���|h?�7 V�����a�;)��/Q�o�A��K�[��gh P��SNך��Lhf���	\[q�����m�l����f�	@�һes��8|M���6VI-E���LA��2���?�����e<=��k��	cw!6���2:so�j�j��=FL�������/���GM��J&��Ll�̀�g��~��t]�Ә?�Y��by��/�n���|t�z�ߣ��^�HPi&����n�c�=K��v/M|�H��+s���9��xԈÑ�87���{��n,v�4�(D�c��*��2��4�F�c�ֹ�M�ϋJ�ѱ�5�vZL�{���G�G��0�9|[iX;Ǎ�:P�3�U���(K&�H�F��M�:c]<.�G;����~l ��A�	$'m�����q���#��9�)���G;��a&0����{�P���t�<w�Zk x�3X�i�&)��%y?V�� &ʺ�[Za'p0��&WTܽȆ���>��fMK�7��mQ���I�YTo�߱:ɧ�d�q[��q$ĪJ��v=�d�A�T�(�����D��"M�V�49����-< �Hdj����5�#��T�����%��ս��?�n���xB��F�>Ef�H�_>�\3�FL��$��(4���rq�eP���{<�������#Ǚ$�R��XC�j�C���{���**L3����ұM@��2�c��@Q� ��z�rC���p���"�����	�RF��;[P����b��u�N��0RV]܇�Uv�:[��!��V�IH3��\;i���v4�Al�����T)��0(��n��.����4q����-k|�,LE����k��>?������r�nٯl�����Z�ծ2��hM\���\����}�~MPI:�-��q)$rnL#k7�N$��ox���e�]��������9&k��M��@�(��M�V�s�Av�E'�~褑o#_�I7cL�I��ɮ;6c��v6�L���Q��#c�$j���8"�2�W�tִm}	����Z�pCǱVb�v�CK@�ڧ`�I:��Ϗ����4�pJj
����ׁ�j؜_����y����>�bb��rmm�<�D�
5R�a�Oi���54���	�a8*evҙ=_m8�{��8��E�F[��!`8�����|�_�t"�?����?�N�O��+����!���G�˶S�4U�[]8���Arj�m��"�-1<l*���s�a&��_Ƙ��rGY�O��uI̪mZHbv����՚x)�oq,�{�(�F`�Q����{X�h��#��霓��]e�س�kq�����MDMKJ=!/%�E�����O��#g+�w�Yڲ�[�~�^V���?����]˘�\�Ek�
�p%������n��B�X�`�ঌ����jI3�N�Մ�.��K[c˖�<x;���O��{�mh�p�A�f+.o�X�`��zR�X�"��t�$v/����P� �e-��IŤ�ŭ:��j�b�y��Zk�pf�V�v~S��V�T`�x�n�S���*�/���_o�6�����X�S��V�Q���Km.\����D���U�z�W����{�͗yή�;�|3E��]�h4u:�[�����^a*d�?�s-��x	ً$���	���z֯�ɉ�bc(���(����Ý{)�l(���L�:p۔���`���߷�a9��*p��yZ~J{��L�O�^"�_f�v����D̿���?
M�6��Og�՝3k�0㒹EHvG�V�OHx��bH��D���Ĝ��%��<��QR�56N�6�|W*��A��\�O�`ye�A��V����<�pT��l�@t�����֙����$!��տ�G�E�$�$�t�����L���v�<&x��"��+͘vb�s)̂� ��/�Vj��l���:�4{�֦ 9lz��Rk�f��-���d�g%d~,iZa�U�=�aw+PZ��À��.�W�g��'�_ai���	��Ϩ��yZ3��k�A���~�OTq�����MW���{yO>�h���̱�U�ū{h�TA��˻�
�Uߊv��K�ss5���ͥP��4���R�A�ǖ�jNr���u��ǅ�]��S�t�(Iw���m��o��q��]t@'���ȇ����eq�
���k.�߆_���S�;�$�>��
X�8�Bl\=�~+K��asssK3�+��g#��a;������\hs�*D�+P͞����G|ϵ2��'/��%�O����M�>�PX�\0[�R�4��dz�6��\A�y����r�q�Ga�&��^ȥ�ˏ/�(��JѼ��&@ZVz�A�Q&Y����VU��fןB�� î!^�A�u�.��/��0D]p䬁�婢͙y�>%76�Uv��A��%�	Q��C��U� �,+R}�L�ZCEH+7��M�:���FuU�Z��85^d�Z�F��v�QId��#W��۟c�!{8B׊���� b^�Iq��	�r�ُ��z��qQ1έ��O�G�{r�Z�kY1�U+G���Ʃz��0�g�UF�p��A.f;ߓ����I�cK�o�_�"[e��=?{�:3I�n���T)脉y�S��t7���5%"M��~2O+�F�	�����-:b�xiؖ1Wt��?rpq��U�(' �+���c>)��,=�ā�4@�}���nEl�+�Du�Z˷���Y/xR�+�ʘa�&��iV뀿OY#cE�}���D�;/ ����Ye�^DeD�B�o	߱�� �u��uZ�y"�͘�� �xɟ�����5�'Ca�gp��§�4�}
�L9GD�c�q�ߙ�H��^N�\��Y%m��d��W)���մ��{�Hg_�Ӑj��r��3�N�2+.B&Z��f�$\ �6��?t�s�>�"X[bje�"�<���SQA���R��ta�I�6��%���5L�JB��x�2����%�u��-J# �̰��;���Қ�y�d�E���¥��<1ә�a��YwY®�n�D�ڣ���<a�D34����.u^C����CH;u��K��ზ��y���.�E`�]iq(/�n�����@p�Mj�wA���_W|�
	ŭ�Uc[m;~�3����������#��}����W�B�}��:X��0�����\;�۬�����U�N�Y��i"��xDR\��~�/ax!v�8c��+0���&
i
�w�L�5at��N>R,�0�9��u�h��kb����x����V�k��4������ݐAz��w��'��}���b���� ��TZ7*<��Z���D!�����}�S^%) ��fimP1e��k6��[���%h�
���Π�`�oE>̑]/����R���Ϫ^���w@�P���\3��iW��7Djy��v�Bv/�i��o ���@�9_�G�R*^�\�[�R��}ȃ�3���Á�Qr+�N���d#X:q��Zg����K��6R�Y�Q^��70p�H<|s�#u $��}K���H&1���b]�\5��j���K�a����[�|�e����VXJ�l/Ď�i[�ό��Y�aD�3�!���[+q��e���/Zm�a��<�T6P��&�i
�7x]��%Y�0�B]O��{}���=c,2�P^�lVC�ڏ��sؼ�b�At�%c$wb~���UuB#�ٳ6��"���� �XƊg2�OA���b�/ ZR�l�L`�H��H�v�O^��n��U颶48��9�ww��,�G��0&R2w��D�5���F��-��n�[;
�IS0(�p�w��P�=���]��^�7�@�ec�����)YF�%�5tc:SQ��g1"��9�H�|J���v�D�*n�=��#���}��ﻨ�� ��	r;���x��KA��xRϸQh{�����a��3H7�6�V����T�:��	��|�;��=r��y{j�m���N�x����U�t��_
���Y�2P��.���0��k���⍘A��]�tU)|����&��mYT���o=�l�+�@�^6#�aV��8!kq�{�m� �g����.�Wڙ''6�
�C8a��w�|(�N�fQ|F���$omucʓ��2T��M�b_'%E�&j�%욌�#�	�y�M���m)v�J9�sz�At"�U�L���`��k˩!9�M�4+`c�Y�����W����
��Q/Y�|�j�q�����Ȱ�¿ۛ��Q�5Z)��=ʓ��z�	u�lώ��>��>ޱf~$�K����s0j��,�.�{���@�`]/���(����˒�0ٺ��w#eUc�9�%�_���(�8����\�Zfik�3@�,7m�ZE	Z�˪���s��a`�ų*�Y��&���ݎ��9a���1��N�G[��A�/}ז~;c���q�BO�Z閞�/�����7�O�cS�ʕ�w(����NT0�ud���i"������P�:4��d���v'̬�z7~�N�����	1d�ҙ��B��˺O*GtW��6@Cգ%WO"J7� ��f��Z05ΰ�}~"�6�����l_�Ն�r ���0�(�ľ�W��f� �\Q��*d�\�
�GH���8���4J���o�kCru�0Y}N�� ���F���W�|��\��+��.��^�>pm�f�:]{�_m[�x��	��K��`Ic&�V����w�Y���m5�Z����h��}y�7"�iW�l�@�C
?�0W�����c�XBſ��4���s�0��:�!=Nٳ*�'���Ӿ��,Sw�M=d1�"���ʏu�ZH�8La��*f�>��*�7�S��fZ�[�)��*���È(�R�:��m%#�$gk��d1t3�h	Gd[�A����le�L�4���W|�����^�.g��p���~��ٱ�Ù�SH�η�1l��@��J� ����e��"�5��"��0��"�𨜷:P���F��A�4󰟷W.B�����u������Ŗ%#��+г�ɺ�D�
�G9���2s�X����չ7��L@�El���5ё����$=����$�3uK<Ք��|` ��5�r�ď�\�nc���gC�%���だ�ePڠ�uN���'�fᖏK�]��ָU�iĨ��=G���rD!�?Eux�*ߞW�ϵ��Ht�����'	{Xu�PYI�ݫ���P����O2��f�u:)`�� �M��ٰg���e
�(o�(p����);G5�"Q���lQn��>��X�*�z�+�4`d�'��;5�V��00S��u�/�yaA�Gɢzr�7f��CV�{�	1;�O��=�2_�����@D5N��l�KsR���U`��	p���I�^ȴ��>�Qwm� I}2�q����>��)����`���KGc�C����$ᘇ���O��'���fR��?Y����R��GT�����v����M�~A�>Zۍ�o�m��F���� ��cc����8x������;�/���O*�D��;W�],S7q!�P�9����,�^Xk!GN��ǎ�L��
1�"L~bH��8WLʹ�m���x�PuoU\����z]D�+��i�@(^`|��~+T�\N.o�e~�+���G^�F�6�ܭv �Y��7�đ����9;	o7��5��7R��a����W���NK�yr.	��+�%D��-HW_��ZC2���4��$:Kj����=q
a���l���+����	Twpri?BS-��=��h���fՔ2q6�vJTn����O�?�6�#P�{]��>��1�^��*�����.�}�-	o���H�^(�A2}_܈�16>�K\7ɷ�c�0�����|m(�b���2��yx�\A�DIa����@ocI6o���@S�)#��x�)Op��fM��pU�Jͭ����=d�b���=�j��X��M���z�4<�������q7�^����6	+�n܇M4d~ 9��悒��ĸr-yG����k1"i���]�����S^������CB��r��*,�`����ӱl;�'�g61����*R��p΁�$�}�����Jc{�@=� T'���Ռek��W4g��?�H������	?���X�l�1g�X���:�v$H�� ��;]�J�M��|�ϔ"�����9�Ϣ$lyJi��k|j�$�r�,BL��Ri唗��)Ӎ��L vz2�_����n���N�;��,���<k��I[����I�Aa*�J8Ш����� A-5"���,�f&�a������6���/l2��b7U M��\֎9�j��ˊA%�|�3��!���n�ux�n|���$�
]T�_����
}	�G����������j�
����2�0.c���L��|'H& 
w�6NkXRx�*�~c+:2G!-�@�k͗M�Z7bH�O۟."[���B�=D=n���洓��B7�Ow)©K����1hX���U�B���x������X�P��7�s3y��G7�lC��������>&<�WR{՝JU�6��W�-� ���F������J�z�`�>��h�<��Ӗ_y�K6�=L�'f�_��*{�hq���8�� ��޿���נ�0��q"'7{�H,�1[�������o��kQ�8�@<Ę�y&���cbrH�a����\�a��/�;������4B��h�B!;�r�B�}gR.�F�F��������Vv�>Ӣ^K�pk(tw����Mp���֬xKo+�-�E@�~���7��wdD�r�z���m�^�fǆ������R2d����I�d�c��֦�N2�z��#�/�K��~{�N$hۈ���SU���Ԓ\f,�m�%]�9գ��:z�`�O�L~���`������b��+��[ ���x���)�	A�����V������P�/�L�E��o^;��#H�f��9'En0C�}���Xc���'_���b��X�s>l��`��5D�_�Kћu;tXF����p��HT�oL����ys��롳�"�����i���O�oE%�Z�q������5�2j�?Cr��!���n�?k�G
��!����;��K�β��} |I��%m�`\	��d��<�!H���]�
�Df��|2�\	.�g9��0��LD��8*1��|pPs���g(����`�ϠM�k�?�Ӂ��e75i���y�?��s����FkSW)qD��s��{hCA���l3Oq�����W��R��`��b�g�%t8ې�6�!A�a2�Os}S$��4֓q��}�_`ҋ�?M+��Oo�f{19����Q/5���"���er�%5�	�N*��Y��ܦ��#qV0��LC\jֺ����=��u��R�*�~ʼ��3�϶��4���6����G� ?� ��3Q�8�J�w���-^�'���'��`L�x��ѲT5�H�9̝f�W��g����l�k`?9��vnM}4�U��ۓ�-�Ӊ�2���I[Kp�{V�i��jAJ��
�Ѫ�v��D"�����$����Z����CyYd���JRs�����72O�l}	���HY]u<u�����_�:�3+Yq�J�^ꖁ�YY��u�e/o�a��22�}ܛ���}��ؤ�c�T�1e��@��I�x%�K�밸Y����e�> �$7XW�GR��W�MG+/}&�Ț�ڑ]@���'�K� ��9���C�W Q���Jiԥ��o��8���y�#�ݯ5����J� U�
�SY�tzP��9:���$�N��ޒ�lU#�=Z�����kU__��	i�f����n>�����n�r��VL�D�u�G��E�R�$���^�xv�UsKG_<)@J�͸_	��~\֚3���6 �óM���R ��Q>w���&k���Zv,F�I+M�i��	�>I��7w? ���e�����=���� �~D�b�H=��r�P�͂�@��Z-��T@>�;��5��w+v:�,�Ձxf�f��ޝ;�0=��[�1#��]q!�����k���WR��G��j��'���ˈ(�z��Q[xF)��}���b��������.�����Q\y�@���5�;:�����Ś��^��>HD�������a��P�X�)�O���쉳#!%bSާ����ho$�w%w�D�9�=�Էj^���]"(�hN8�w�l+��Z�N#jLW� ?�[pd���/��9֨C�K�|%���� H]O1�i��T�a���
Vc�+t��_��f~|��Q�
O��@���M��"���=�fi�˻��d�&#�3���,R�{�,j+��P,PiuM�j�.V��
�,9�2v�ppoK��|h~u��T>q���	���_�=I����[���#Yk=��������_yCQ|;�,B����Y��^�*A*�CYRY�8D�u^����#p�y/ �Pd �f��GW[����6!K[g���m�y�5Z1���$.���ם#û�4@�[��_�ܚ�'"�/RHg�� �<��e �����z��ɭ'`�������mA�z��	��[����$[LZSMjM� �#�D�!ê��䗎Y�l�3�%�@�2�=�:؊q�ӎUE9�4�إ��e�Y�|$�3�HG�3����m)��vGoށ�@�LEW�z�@G���߅(����`ط�#�+�Ԃ+Jɲ�$�������p��	��5��s��0�R��rh֫<���>�24��?ç��6�/��qS���a����\V���m��-1��!�@�>&��ZJۇ��.S	5+^�`'O��f�NЈv���5-*1,cR/s/�����=!D)XwBG4IijH��*��6ɖ��VF�p�����#'��2L�~z��E�Y�á��(�R�@���� �mC���bF`B��<�\3�i���*5u��ȑ0�-#�e���*��O�@�q	���#uۻ���a]� �.�ˡƲG\�v�\B����b���'+�q��&�a}��<R�Jutw~�}�
�2�}��1�b>�.�sY�W�]����R��-B�*�����z��2>����F���wn&��G=C|[}�;V�q���X��\�՝./Q��ScO�����~0\��G�C议�\�\��k��BE��!�D�1k!���Pb2
��AA�_�rH;n4f��[8&��}�օM���"�+����.M�7*���24n@����l��3�$���x��3��|�Oq0�jW.�?)� (5� �ٜ��jG�R	e�m��I:�SF�S�u!��\��*i
���ٶ�Ĕ���o�g.�iץ�ۺ���W/4���wM�xɻ�����m����!�2�^�TG$5~�{�j���K��9T������V7r�-���5��@��w�g���z��7L�]�-ʓPbGFw�oQpsI�%$��i��lt��5�k����%Kѣ���h��߀C0q��5�,�f��Ҥ�Rw�.��� $G,(�L"z�x�b�P5ŕq���OS�uޮp��M�o�I�K��.���)��X�nv�l�%NI�r$e/uuĤi��f6s�V1������^�^6Nآ�u�V�:M� ��43iS�;��YU���"�m�|M�:2Е��������"U��]�+�U�b6oS��j@�^�z�]ٳv��)��2\��3lc�n���=����<�kC �4����!��2`96C�l_��������qɓܦ��=�}K�I����,W�5��p���`�5����� wg?0��E>|>���u?�忚P;#|��9���}��ն�U����H�!	Hq���5���H�� *t����1S����r8�l���R��\��9�V���2Ii<���~E1�;��RZ��!�">���s��翖��U�}����;�@o�<d��.B�x%�������c��8�<�6���ߩ��ߪ���UЉ9�0DE�����J��,
zn�-Jym��pI>�F��OF�M�"�%{�D`J�mc�&����Pr�5�7�J���r���2e`���E���/ ��듆N�Bo9��bW`���):w!뮰�e�U{y���ݕ�ף�k��V��Li�p��g����;}&oP/�[VU�u�Ψ��i�vܺ=�}Nk-f��a�-Eerɮ&�G.`C���vo��m]/�[5P�R��uwDLz@�ZJ�.[�q�#m���j�&+S2�H��q�bt��8��Wސ�;�U���4ƀh���Μ� �Kp�Lʎ
܋�k�L&Q�Q���~�����d�U��h����c������]�Y8�y�b�3�{�'z�����sb�K'�y��YÛ��pàBM�=��h��X�z���G�:Eh���{G_7����t����إ�rÆ(��/���y+��-���{w�W�Öm�fK+��nƤ <��;b��� �;{)��g XPگ!�A�ҟ]�:��A�2�^K�8f�O_��.Y*�o"W�Y��ɶU�w��t�h;�	^��wU�v@M,���ꇪh�g�I�_�]�h�_c�ǁ�-��b��A���=9���"��gY�IL��Y�ۋ�x��|�)���jE���/�d:x�I�R^�-��eśE��-��8�.m	�����|%����^"��J'k� �7�90{-�����g|[L����<,^+�|��7l�j��Z�6��Ԇ1�<���oLe2�B�gd�UE�p1��6�o��ve���ܤ�L�tP+����ϔ�~��	K��1ٱd�ٱ��7q!�Ҙ~��DM�	ađ�>e0o���J	K\���0�p����-�j��@�%G�kW����Z��1Y�2i$��ұ���I��Bg�+	�D�����U��u���2�(�#/�֭0��W;/K|�9G��܄T��O��B>�a8����/o1�ې�:z���1S�X�_����eՅ1@g#��P|�*'I�l���_��V�K3|&�C���{�Qtt,���r/���/0��ǌ�d+|L���g�9��8����F�+���;$iN���k;Z'���4�W#�'�Z6��o�˞�t�-0��nC�+��(D#M�� ��w��`�k�=���y&�S{6s'�FY��������	�'�x\�V�Z���"��눅&w;��s�`G}�0��n�75�I�fvonCI�˞�a��PJ!��Födz����Ge3�ш-�5p5I[A�Bp��`*l>	�aߌф�~���'ξ��u�2ڿc��ް�3�y�Y.���+P�d��.�%`m�ɿ���Ho:i)��y!����h�1��S춖��m�3*V�*O	�sA v{��t�e�S֐C�HxW��:��yM�u������"NAV�>QK��ҕ�z�r	25c�Laf��PvY�ӎe^�!�#�E�l�P����FK��	`գ�w�ͱO�N���u�R{�3y���%*)^�ס�-Xp+Vs���%	i�2K��*��_���u��u�;G�1C=S?I����z�N^O��{޺O���������-N���^U�E�0���矪VĤ;���y�AM�7SdG�&�	vI�^�y@����^�{HtK�?�r=?ǩ7��Vb���mxEWG�da"q��>��:���V�D���KQ��@u$ �J���L�c����v�����Eҵ�ƇwH�����D驠�D"�u��s�#���o��m���q�EP@���q���b�(���NY�G��jv��JN��U]�x{�������8�����4-���xh'V���1�e.�;ڥDQ�w�A���!�����(�븊DX�w����i�q��EU!�9��m²s���!c�$��gC�av���8t��t��e�:O0��MFKǗs �``rnE�B�iH�J.����o!;M[�!I�p�92��'����(�G�˳���F_��Ϸ��TlJ�=�~�a�"H��\����{�aϐ�y٭�q�K*T㭧�@c�-Q���͙V\0L�]��+Ӓ�-so琝��E���
e�k~�`I�uhg5CU�%�	��C/�>��y=5�/����:c+�D�|_/���)�����z�[�x�1�`��3�� -K��?C��b�dZ�\'!\y����x_��̫��I!O���8���E̩iy.�oFZjU���[B�96��e�Ү�Y�;��2��Y��H���$���:et�FW�/!�)����w�6����:��!{Ƀ�X��^��o���O'ak�:,�*K�+Eb�4]�Na�Z�_^	|�r��0Q|���[���I�R MZwر��YHo\�`��v�Y۔ݝ���"�F����B���
gN�^�i��oSǼi�	t��2ybr0�g����Q����J#)�� �\�ٜN�Q�.�P*]���y�}�ǳ/��O"�Ϟ�K�X���,8QE���p�J;�@�%@m8R�N*>!�=CYM��0Mm�*F�zM����KD��m�h�$��������ǓJ,�]�� Hv� ��t�Vέ< j��)���������z
}R��H�|���ƜΞ�JdBu�Op�V��BaӴ��������'�rk��-�RcFw���!���ޫ I�p	_�j�4��9�H�w�tۀ�=��r5��-�?-VJV>���{l�}L#��1�� Mo 
����J$��'���^6�ZӍ�����Z�1J���q9'"�Ca��]����H�UUȪz�׫9�f�p���S�D����y�[jIF��N�����@_4�S+A��z�D�yRag+���4��'A]V'?Z"�&�W����+��i��@r���:(�D���2cz-�}.mO�3+��y��;�#�Cƞ�n���N5�D�q묐��--ށ�%mk�z��<_�,��>i�q�>n�l�Eu�D��o���ta(g�£S�o���=,�>� ���S��ě�3��4��a�T�KX���.�?�����Z�i�����S/j�ɥt�.o�%�ҡ��}�s�kB"�glk!���5j{�P��5BBJ��xʤ����b픈N��? m�5j-�̦���������Ȥt�9<*�w�5��ٌ�[�]u�`��R�l��L/�	3����/��"�����y�`I���_����k�j��Ƒ�O� +�
���q|�Ja��[E�hZf�.�$�&?7l��!/v�H>�-�߉{bH�������Y۹�ul玾�g��Ҫ����!�`�����X��*2z�v(�7�uzp!E��4�=[YiH7�*�8�c���C�e�S��v�.�:ST��������T�Z��@rC�����_诐Nh��{U	�.Hi����=�� ��:��2F߉���f�����of����n�ˉ����4I�@���i�@4�l3�¬�7����u���V�{5T^B�Ւ�"����D��:,X�l���B�nƮ5 9�m=��Z��^R$����\�9��VO�#"�	��I�XDK�Pwbn�JE̡@*�sD�Э�E�Km�JY���h��Q���X�����r���h%\B���ٓ��Ϊ��\!������.k��6�}���v���շ-�]���k'�޹�~�e&'��G��h�!�;=%j��k���~D����vJM�"�T$�lq� v6DL������jA�d,��L�c�!S��w	E7�F��2�W�����hh�g`�O�G��x�w���*FS�O���2\�GS6��tG�� �S^$�A��HG�>N�ɏ{8��9��б��]Z�8�|ѯ�qjT��W��P%iǻ0��A��K��T]AC@��P�V���8��s	G��K��FY�`46W��;i�̝��*Z�a����Q����B8O�P�nk�B|�y��s���2�@��8{�Ϳ=�|�(J�*���I���
ti��w��ħ�X�KV��l�/�4C�6<�n{iu�^��Ӹ4c]���t���_�4�2d���bd�ivI�/�7Ȉ��@�i�)wW�q��ޅΒ�����g�1�K����6� ����W�O��'t��jW�-2�Q��T�|�$1�є��ׄ�u:"�Ъ� ^u-1z��j2��=��	�x)�l�P 3�!�g{L)�Տ�ƶ���OIj�A-gZ`U;s��ЀT�ni�)�
���-*��E�{������/q�d�/|Mrw��*e��_�3�� (�l	)y����;�[��M�=Q��K,�@��:�?q'3�[wiKrµ_Xi&�vUfΏ/&��0�Z��c��h�iH�\a�f`<�C���&�����dp9ً�z\�Q��OH����O<=<����3��w�֠f���˪���u߉I	��"�L�&�>s�� �i�MqvW�_��>)"HQ�4��9�G�Q�Ջ2y�G��E�(��7�n��T�G"����,ۜL�D\��a;}�}�Y�WlǷaC;+7��+;KJ���B�B	����!�Ч���C�_�
_]�����q�i2C����>���$ v ���^wER�;��B��to�E��;Wm�m�(�#Ѭ�t�Z��{�{Lnn7F�hK7���iO��?���l��)=�r;?�/�t������De��W*�{�s�7s_�ɧ�ez�h��/ZHkgG�����XN��3�J�p��pC�`��E�D`�mG�������5;�	P��;�u��(�}3'\q�U���.ǆ#���?J��b���Ɲ�D��y=����}�vƸ���i���3SR��7Վ��/T��4��b F�O�)A�@�H�/�7G�@/��^z��l�����eq�n��"��"8��X���I	tG��]bk���H�~5B��ɞ��d"���Ѽ"l���kx�}���n�*����X-Um(?�,�Գ��5]2�楬����h��"{~��<Q�%�F���&�p#.�J7�P�����$e)���ҙ��HP� �0
甓ׅ��\T� k�4����X�p��Gm�ob��'�j��!'`�ޟ�ŅDs�V��Q(U{���M���h��E��a�]�9������]O�:�>3> |b��j�P`v�;�P�?��T�����A��N�h>1>؊�=�|щ��B����p�bwp�1�i�9�{��� ��hE@n�
z5��Z�L�ă����F�����ݬpY���N�U���M����0�����D�V�YH�܁���]|�s�I�D�������x{��F�<��3��q9����G({�����b��oc���8G 8��@���eY��B�P�O��25l�f���	�6�@�cu�Ñ_���t��Mi���������!���Tx`o��r}�DEQ�X������Ԩ?q�	H��!��m���F'��[k�o�p2��oUZ�(nB�K�|*c���>�s��6����N)Z�ƐfkZ��p���ȟ�8��R. �u[���n���9
��Z4!��<-�"b:�8D���Pw���N�¦�{�9�@�!wv�=	�#W�S�F��DUa ҩ���*Օ��'Vֿ���@�U�a�%H��zl�f<8�2R� ;C"X+�Zb�T �{�1��^
<�-P����J{��Ҡd
<�;��/��F�W�A<mv+�_��16Y�����q��Ѣ�(������a��rSV
7���j/��ca��ˢ��h%����q,���l��S�%�o�`I�ŗc킬6�vT�`.��1�����0��j�x�n�U��������0~@F{�hm���خڿ���oR��Qg��2���p��ǃ�cN'���}BLA%���"f�0����X��n���⌶�XR�B�ǭ�u�Du<�1�d��������P�zSP��R�RNN@O��D�[��? 7���`~@!�+mOu�Ƭ`�S�*�`����}d���
�hc�J�B�C��8���+	,`(ɠ�j'��z�\��[�K�+³_��j�z���M�,�o�%�AW�m�\����ԶkH0�R�j�/[$��,,^=�%|��8� ��W�+�ʹz�<�S�a��|�{y\>s��mK��1��b?gU5mG�?�j��A�� ;�S�}�}�J� $�Қ�>���eCdѡsX61zj���f�ڻ)q��]��|��'|��#�ç�I;>��KZ_%����VJ���\ EM$EĶZ�;F�`@7�2�F�~��;��#f��EI��N��c���n*��i��kFg<�������5Y5�&��!v8$���Q�dTTF�y��68�L�y1�q�v^}T)@��v!Z�M���"����� ����n��(�)d���I�)� ��f����Q���-�ډ�I}&7���G=Y��z]bxt�� }\�~~��zr	���Pm�����2�fk�
W�Ը���C#T=�n ��<�����cTҴ�Ā����;s�\Q|�K{�|$ٚ�)zr�E��L��~V��)Ǣ73>�P�Y�ľ�����8��	�L�6-� s���X�ZT�v�����aI��ndG~w�J�#����M~x�q���Ӣ���LZ�o���E�~Ȧ�Z����,+8�`ί�:%xO8��G����!�vhz�rI�K�6���=�7��jS�x6�Yo��^����y�ݳ�<��z(E�9��>��<Ꚑ�7���o!��>EP֛nBҙ��v�9�}�̓}�k��Y`|���\���p�,�Ѿ| ~� '��/xj�hp-`��_���Vw�h��|K"��l�.y��Y��o��f���P�	�U���;,���z����(C��Ix�Pk�!�&���Y�t�D���Y���@~����}�����^�,�u�C�(f{�T,�����#�{�Fo���;ȳ��&�����6+�i^�w%��m��΁��EGV�s�]�T!cW��p���W�J�����������_����-���ߐ���������|��]U�hĞ=��*]w%�
��(W=�b�D@Yj�Q��/|��R��C�X�I���:}�51n2,���S!���s��|d v���#y6SS7Ǌ�sd	�\����q5gl��1�vI�4�)�ٰe�@���y}��t��xuߩu	�P��n�:����\�۰9�6��j7h|�.���H�!�^�=/�hB0�k�M(�,����&*��Q��ߓ�o��'���	-i�NߞT���9.�����u��g�Xf��}O�GZ@�)�
�θ҄x�h��Dx��s����Oo���u�=v��Q��Aʼ��,p-��3t@�jd!$Ȫu\�7Y:h%S: ]��2*�:��{����e�������*[>�r��Y g��������=K��R���:Y-b�M�s���y��L]!���sJ=��nS{7�m��� pŀX�Y����?uto󻪪�I�	'!�b����j6.1�{�2{9��-M@��C�z��a�p�G�S��[�(��0�*��W�C�[A�*�'��
pA����>��>un�����w��^;���O�e��^����W�"�E[�؀~ g�j�n(h8���ȩp̷@�>�7�A�Q�
P��ECu1e�~�o��Dswĩ#��b��u�g ]Q^�"v8�hfviV�]�
5(��ֶ��-��_A`$����&U�#�����8s�#�O1Ð��\
�r,�!��M�`L*��8+��A\�����EJ�룆d2fs��1��&YM�9��)����"�c����B9AU=��7��-�5 ���p�Zn����m���=����a�ۉ�w��x`����:`��³l�咄��w��2��v�?����4��tC��$����v�s����o:����2�U&רƶ'��~��ez���
\Y���6 J��*���)E`8M�f���ݲ:
�����EoĢ0R�*Wنd`V�o�˖<F�T�"�D�L~�L@��K�f���B1��:r����E�!�?@M��z:F�p/�YxӴ�j������v��d�BaC_�*?�~Z�}T�Cr
[֘
�q��/��(3�WC����Z{�91�[О9��eF[,Zj��|;�R�Aa_�K����,�(��R���'��;�mxf���ly|y����C)�(�઱�66�\���q2�l/�v�I�\�j<uLxq�@�<�mC��ĕ�A�FQx�����r%�J�(�LV\R �h�)���X��-9e�)*B���'FW�W�����+$�~�{��ʩ@G�v��S?>X��0ȱ�������V��x�`�hOo��%X�#��4!C�aG~i�-������|���N>�x0z�(%�ZJ�clK���&��43\�ڭ�ZoP6K���h��6��"��v��R�8�V?{�7ŏ	;ѵ���}/��8	�~�9;��n���ߡ9�������`;�In��;��V���N��a�7b��q:�$�@��=ȾXs^p��V��l�RX�}	��}yWF�Ә�� ���#<����>�B�ϔ�'�UM,��23�0�#�}�����!f=T��.i���q���)��׹k��;d`�0��u��ϵ[�v����ӭb�S|X��Ș�n ���xHJ���{�G��~�J[w1����(�e�a{�)�m��l:�5�|���	�Fػ����5S�p)��Ä�h��6�#�z�}����M%Pe�B���/�������=�Mk=��E&\�_G�t���Q������� ~���	hQ��B%���.�#����u��v�����6�����'�$�|D��Uibgo�8��m�`5�kG���&n�5q�v��oP��p����}
B\N��ͽ46�L��E�NO�@s��Ei�����47���3f\Z��9gw1%E�0&�U��x�:�
���mJ����V`8�*f�'U�����_Ra��q4�њj�srz���l����vDO���4}pe
Q�����]����9��M������C�oȣ��~�<�.fUn���7mT�ȉ�M��{�q�~-���: MO�N��H526��ԩ;s�щ��"pƺ��z�����s�Y`;�����c�����3ƽ�Z��jD�'�[ѡ�	Jc�W�#)<�v�YS�ņ\n�d4����SG�7�5dQ�$��=�Z�������h���\D?���|�1L^ǘ�^E��>�9�M��+�0B7>Z��_�����8�P;���g�ߒ��-���Ȗ>?�U���헭��wԃC�o�?2]���O��	^_{3?�`��:��DT��=�k8_��!n$%I}R�'��s��B���Ip����@�;_e�{��G<���KG��p�W'z�tI��� Jh�a�����βK���v�b� ��3-�-Z�O��V7pe�qZH�R�dc(ׯ�r�(-4A��K�F|�.�}'}��R�߫���������^mLL|D2'Q��FY8�Kw.�����z�X�|s7�(�C����¹�SR����_%��Q�զ�t�<0X;���A�9u�C����e3CTN5Α��YhR��C�|J�6��B���Ĵ�O�Pn�M	������F�o��g��5�s ��]P}7bV\5�[�<�BjB�9�z)M��`X�x�̂��Aʭ�iv�a92�p�R���>#��F��g�������vmQ��|X;��fD/���$ {+�6a ��71A��yx��bfrM��O.-�a42�����Ԑ�|�ʞn�aL %8�����LC+� !��\��|�������bb���)\��3[��F�G=��(����/�� �d(���>�U�C�P��>��Y@ �K(�B_�ȼ#[W-��p8B' /�w7��~�	q]�ʘ�N7�ҟ!q��M������9��w����8d<� lP�J���G�=��*���ؓ��$�_O�R�x�|"I�nt�ԇF4���u}u	��")⠋����6����?��iRB�G��|��g+��Rԕ��~{�Y����]��������.*��s��H��3	�(X�V�	m~�#I�����O�o�W.�v8OA��ER�\(J���s������1���w��	���=1�s#�XJ)M�;{+��eh=�?u��s@�FY����A��e�-���'���z��Qh�_J��p�'.��yw+
���7�y�Q��y�6Ӫ@�_sy~�X�i�����|���i�h�����#��R���`�N���k�F���^5�?�h���SEO*��J��s����� �6&)u,pS�,��W��Uc��Iu�,��r�9�C�f���u�(n~�2aV�)H-�9�p`H�`���v�6N�����b����5�c��㆕�Qf-��v��Y��g�.ދ{ʆ ��f��n�5�f#ϑ��E{'oRr�d����r�n��6᪩���֑��hۏs7z��)���l�(ܝ7n�'�H��+��� K�T�(2���;��ʺ��2
$~%u��Ĵ���NC�o�lӳ�V�#V��I2�Kb�тF)	˥[�3��^'+��CHh��C%O���Zū�z�T"���͝�X�QJ���� Tx�)GU���l�!�];�s��&5�P���C�\�������;��ƾ�}RQ<ysjn�*���������`��"�a話0F�Xh�=K�<�-紴�Fx��v�^�XCĜ�Z1�^|x����xT��}����c]��ڲ���k��3fQ�9�#����wE'��Rt��#A���`�i��>�g�����p�����F�dYz%S}��H���	��3�t�&�3r�$���_�x+@��J��y[�E�8���=�?��Nr�t��Y�c�2���)�Á_U��q�0I!,E��r�U�z5E�}8[./i���o�~�,�k;�sL��H�%�v��6y��h�Z��Ȯ��'�9g�[���!.��v��#�;`�^Gt/���/SU	@�Q�/d�6���ܝ1�R�:"��p;�1���
\�ϑ��䑶0��������l��Q��Tr��$�׫��$�h��x�!'�#��{�'3��H��� !cc�"-�A�u"V�Y�y��K5���G���-�2�����@ �V�i��˱k8}�D�糊GH֠_�,���t�8`fR!Ά�C���Pz@7;�����6+u�D������g�0W\
����}L�Qm���mc�&)K#SJR��a<r�d!�\��YB�S=��\.�rL�yLy_]E3h�N��<�P.^@�(2A��On2	�	�V�`�`�F�z-���Be�$�ٺ�x:�W@:�_��D˂%:§+{5��4��� �b��z)o3�uh����1���i������S�7�v.;o)^����Y
��n�Ǿ�պ��#폑��c�j����؆ꠖ��-�7�e4F(���0X���O-�Q�:����%�P��dz1~U�L��ݯ\��9�/��P�P=�A2��H��9s��o���X��!���O7�n�Ǒ-?���ǚ\�uG4�|���	��� �|�d<f'Al�\�^�E�m�[���c�i�xA*�IP��W�@l�ԟр*_>{���S��\��6�K�>j��Ì2��Ӭ�W�%l��,��C���EX����C�!=h�Ls���ˡ�������Z�.ϳ�=���</���n��B���v`�W�]U��_c����������w�9�i���F��-��ֲ�֣#8`�n�XП$+��Z��^�D��N4K�Ft_�r�|/���Ja�)�O�}�8f`��!� ��!���'U�7���	�1y�م͞
�>�i�U�c��� �U��[~UѣG\�Z�H>��V��;�V�@ȸ�$d���%�P��w�M
ۦ ����w���o�P�W���T�I��*:
�$Y-��2���H5���q��7���_ך����rC6����~�H�ʜ�h���[�fq#vT(Y|X��[�xXW��\�H�v3�����;��b��5m�QG�����GV�I���v���-��"*�核T�y�HQ^��O.x\��%<�{�h/X��2�e��ȯ	������K #���ڝ8�\HZ�p�t�y��Ja�:�q��Ed����[=S{Y%�H����4�h�W����FlF�#+��SfQ�SEZ�8�����=JM�����7>SW.XsA�QKYV�\�Q �!��Cf8 ��#�P�b�r��%F������C����B��B��|��e����RT�r;M�J������=<��!6g!8��IE~�ϛ��r���q��A�d�-���4S�ێ��qm�N4��yڴD%�4���%>e���g#�m���