��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)��<�=�!�hF�|��!�$կ�!
����Ҍ�&ј+6;��;�}Ȇ*�Qǲ78|��g��g�ɾ�>p����nG铛�OɊ�(�3��\
�Mif���#>��4����C����(�}�b��?yr1;�/bu˞A�����&�O�g��͙8�R ]@���� X�%k~D�'�EK�F��ݎsM_=��wBd�����v���o����8�[����e�1}�>x����L(SN��NK��R/�e��ώJ�;�c����4���f����V�+rC�:�꯫� �k�7�\�Rl4N�~a�x���ֽ�?�$���ϓcK76�=��`�4�o���e|���q�N;�!y2�\y���0J��맗�kJ�20v�~�&�[�r��&�)ipm�5Sw"�4(�|��ϲ�Ub׮��)��r� f�Q�� �hI$�2����~�q+��y䞑�I��b �-��u��jʌ(Bn`�����<#Μ&]�FE&u	ʛ��٪	=;����y���_�m�{[�r*��X8�c���M�T;b��s����v�=&��+�Ԛ����1`�L�t�P�������%��r��+�娒��u�!��[d�G��K`,	ѱӼ�F��~����N�Ŀ��HǊ]�RG@m�Z�����0v��0v������}����,�rQY���Mj��v~(9�ΜC�zn���#�s��kܕ�=�h���}T鍫n }���5)eKH��%B�,q���1r�)�;�>�7%!��6��A˭��x�mV��[t�#+9��}D�~0?��8�ff�M���1Ԓ��G�����1����pBGaB�ߘ� V�x����n�s/4���K
�0�Y��*���P�5��>�H��m�3��}Z��҄��RP�r��Fs�꠰�n���'��	��;�	'�V�G8��ӥ�)�a����19.3_h��q�N��z�/�W�d/�6쇅��a�#W��_��QJ Q�A��1�������^}pB�'sU-,�V��Y'�2��,m�M��NV����B2����˙��r��������%�ZyB�h��7�/�w:��f�e5�
�1x ;��1��d��詻=��_��$Os]/��AڋM���F�	���Q���'m%؆!��5cY�Dsѧ�K��RD��tE�mK�z0��pJ���w�T2���)�G�a�J&佡�K�p�OR�|K<�J�C:i�\2T�H�n�����b��#�_
YZJI'y�:̘���m�;X~�����\�)X{����WN;���͡K�]�J�0����ܬ<�s�PL�*]&�����Vh�~�
�i=>?}\��FCBx ��*�pT2��0�P�t��ݫI�����:Fe��5�U$�:��kN0�qw�tQB��:�b�#�Y�R|p�u����F��=0�N�r����m���u�	�P�;�dH|=+��+���OdA�Y�3g�_�툭NM)2�Y(�����Mt�1?">��+���P��}R~f��Xmmx{��*��$����:�澁|~��$�O���@�0/b^�5L��~�	���n�5_�D:}��Hj\xa�ld>��lyZ��]�d�!��%����2*+���\\�ol�ė�A�W��_��9�T���Ip<��3�u��"'�C�L9�eS�����ZC���X�iRx�u׼��7�I��8�v=9�2�M�[Z���M�Y桥���!���i\|3^�7�l����E��_����Ѽ Z����=1�t�ڌC����8��F�t΀$!]&S�ZӮ�<�S`��c׆"�ΛEH�O�R��b%�p��,�.��TW�JQ1�G<)�?�E�&ʧO���/V�j�U��_�*�W(^k�-��'����|�4��)o�r�X�1
�/�Բ=��_��]�	k�tx��C�*G��� ��l$ͨ�OY��E�7�y��ٯ��B�"A����D�ͷ��j�8��.��3��h�y������5ۊ����VW �f慠�I]� � �zh4s���e͓�\����un9�,��&o1�.�����(�>�����~�?."��r�ɻuR&���XV���n�Lm��'��wT���O�D�����U�����1 Ҁ0e!Rg1�