��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O�u<�9�F�|܇�?g��5�I�h�Qz��w�K1)��t]��p{�u͑~Y��7M�(u�w%p�	��	+�`W[�'L�������4sl�PqD$e.�n	R]a�S�A]9�L�2�f/R��&��.pߙo��o©⨪��RF" �����	�Z؛�W�$��Jm]�g"�|�������(\��w7!���l>'��h
���	�U�7<|��e������*؁�!�0���4Z�� �窐#��,���7׍&�Fm1�BMZ2��A�V���e������ *<jZ´1�c����2v���뭬��߀V�3k`����qDg҄��`��.�M(%k�{�Ї���8j>D�uD����3%xݨ�1�u�(�ܽ�w��I�K�\��/Zo{m�0���YC�	�Ly�]\�\�@y*�Z�~]�����qo<f��ޠ֣d���d+��;a 3��+}pf�SN�|��o����^�0��$�(W	��.>��ɕ8:����{��>p<��	�H#՝����.ߨ�K��M�fvV�7h]'U�U�Nr�[��6�h:�*��H�`�/c$-{;��~��Ķt�$ǝ����eֆ��b���\[���u�L!=����:�9���Y1��ۡ<B�	@����8PvG�E)��$�h�h
_q픃)�.����בP��-i�����%4P�T#"X3��9Z��ocB�|,�b[N��z�����M���t�E�/+$#�G�X/:���_��7�rF��|�蓣.��u���|qVu�؏��5SP���ͤ�J���=�'d׆m9og�>���ɸ�#o&���3���vL�J�U�k}�T+:�a p~|t ��
���o�s�Y@I�&"��ubDS���΂����&�\�s��td�d�y�M���%GXk}�H��!�m��Βjj�9D����={�WXtf��⊘'��2k/��T��c�>���0&<����]5�{I�x��Ō�҄va���]L�D(�ǮVOq���b��2�/4�~�{���wQ�� ":�G�.���1e�`�����O�Y��2���:Q9�.n{�Qbj��+w���H)���d{Ɍ���^l�.�֦,ضuʧ���=Q���T�������<nl �)b��őESL6��t�e���dʰ1/&����!��'�-�db��Y���6-A8Oi��i@�ҕv�6g:�8��B!�)�4�X�|�5�e� ̂B���b���m���*�®�h���5h�F|���$q��#�,��Pݲa�{i�XF2��/� ��s]�9J^��n_=+6bV;?q}���{6��v����3W71e�>I�h��y�<iF���P����{��:��	D!�7��9X�KS�-��K�F*�[�T��&�;�r5*�e�h�z%�u�I�,3CJ��F��wi�*��+���҆�Q�p�*(�]&�[0@���;(�&�Y��۲�81�D� ����=��j���>T@F'�8V��Y��'�Sy�>RJP'��a�Euɝ��籇�܆���pU rd�6���~����7>���G��A)ai��&QA�ǜ?���I���cw2��TfLy�.pH6y�H��D�)WG�k����Ԋ<�O��E��P��h���+L�w���Hh����7��M��g��}�/�����A�f��+/����7i����ˮ�8���D�y�Y�y><iE��To�Z�v /뻗$LV�;O�`IDPG��3��*�(S���s:O9\�T�G<y-3r��� ��-b��C
�����R�E���Z]�蝑n������e��w��Q�X�N���>�d���\��x�B�1r�Sj̇&eg>��ޏT�LN~���4q��<�h[��Oי��DxER��w��q��`{˶E���z�1:{y�xizY1�ĩ�h@��{�	��w�C��0g��_�^���jR��wΧE-�\g�����C�I؏�yrD��w�K%�n�� �N�$"!���J68�[��k�G`*e�2v�]b�.(9��M�V�;:aK��
y1�c��b �g��3'~��רC�RS��$�8z�
F�ӯIӉ祈��锔`~h&*��:�*�Z�yd�"�i*���/s;��j�y�Ykڋ�tT)W`�x$���8/ﺁBT����yG��b��f�AS�۽ ��ʫ#������>�^|4��`��_pظ-����aYb`S��@�$ΙX���u|�w��ݦ|�Z#k��0�v��[����j��Xr�g;�X-v5�D����r��g'���=Ɂ�w�@	<ޑ��M;�g�G�T��'�����_�����"B����W!_S�7���/���ur���������!���Nl��{=҅�7�S���*��">�����?�Q����r��MQ��DRh4)�ʕ�]D�4���U����o��=֗2��|�4��5���O��\0"r�i?2
�( VJ�)<9��ٺK�:ʛd�M�[�w���P�r}S4j���)5g�aY�J�C�e�\S�-ww3�3W�3L�<8�~5Y��O^
��uw�EN�)���V^-2���{Ƌ=C��&�M���h�ʪ�p�~c�?PaT)�@?�с%)Mջ�cH�QC�ՕTr��_"}2~����2��GϓYHkdF���S�yv����/��{�N�)��R/R�Y\{2Rbf�W�����o�W�܊��e!˩��8�ym\��lFu��*�����Pp�p�i>3~у����.r����~����W:��q��>��U�� '	=Z�E��A�C\��er�+�:����d�mE��^Zc��i3�O��6�N��Z���'��ӹ`PL�����S|Ke�P�@߲�����Q�l�yx[��[hk�k�	��%��4u�c��p�vR��[e�v���w���R��� *�7�����/�Y��o�q�,ͽt�����\^s��ð,[��`�w�"^a+��^F�}����\/㬬�xr�̏�̄�?��W��a��^��)Q2��_�|Q�j�0��.�q������'��S8�i�w����V�Z	���)��X �[4ԙ���M,᝙JEa�{�JC�bhU��P䊫v��i��������O�	���n^g��)�ٺ����|d�oTW*ر�YV���C���yMꦧ���Y@I�����sd��!Y�R�ӛ��}�u%���PU����S�L�-����Q�����,b������Q����4rz�F�;c�I.�6�g��%���نNG��y03�M�-�l��]��M�b���+~C|H^� ��v�8z������I�[�0�L�p��)���rNk�e��𾅪����0Z�e��@���{˥!&5[�7��	%#�
c���AC�}���G�1/�}w#d$ &����8����,�L.��_����?��|�z�GcIS���$u�I��SvM�e�������/Kכ�!�)^G/�HH?���y�b㭕<gL�5�Q����8�GTS���� ��LȈ�=���z��R���}��8:`�o��[}�.�6|�zm!��L�)��-����BE��E��)�A�i�Ng�V���%xH�'PY�"�����zr3��~|4��♄��[�и)$X]��i�4t����Ku���� ��R$ӧ@�>HHi�b�D�e�N=���ɖ,0�9���f���]˸����Xh6�Ns����ӎ��n�+� �p�Jy��T�dF�p@���=pXax�1mS_8q8'wf�Hݙ{��{PW9�'�c�I����V�C�$q��҃qo[J�����������������*s�}m�5`2-�K�W�=�!�����"9�)*�	!�e�ʀ�2�z^������*7qG��OZ�c��?�������%��@Bx���c���P\��[i�=t��Q��P��{rn�&��zM�Gl�-��Y������ײ_�����/��Y ��BK{X��$q��>TP-U����H���ܳx��ܰ#zi���@Z$�p�j�	f�wL�ld�5/�`oo�3F���|�ǋv"�*o�h�N��`W�H}8F�N�Ċ��I�{^�h�o�]��z�)����(~z��'�q�=�����g��iG����Dpy�ɝM�#	f(CW�0ފ;�w��ֶ��N(V��������!<
�]~dQ{ϔ%�������5]�|��x9�T����;Is��:i�]s�bF�kS�*�c�1#S\�|k�U�ᖡ���ɯ0K!�j��-$F�3p��~�̪t)��b��:��e��+�\���Nг68����f�+��G
�sq���k͏��,o��|;��:+��?�b'b�;��!�hc�s�:�쫱r�'�>��qj]���[�H�J/��Q*�mйY�t�X�Na�!`e�䖗�C��쏵����M��s��������Q�2�Xo�3D��]<��0k�x����d�[�B����#�^⌢����T�	�)F��R��.�s�I}��=�|g'�����|U3+�(G'H ���E�v�gD����(�T�x��MR,!iz
2�鉅��{-��m���l�lxr��Ϋ�^�#xb��z��ݺ�{��9�03�<pm�#����8�l�C�CДV(ۡDj�>���;Lg'� �x	����r�ԅ��5�7)�KW�Z����|����-��_OQ�ژ���.��q�X2�S2�}��W0 ���C1�͇]v�RJe�ĥs�\�(�:�2o.��3.��?%�n8twH�,y�o'��:>~�����I���>�Jv�n`�3�ܦl!?��{�?�T�FW��Sg���u��� ��5BZ�u�9�`��0��0W����w%�k��Ճ왺�����D�H�g\���d���E�f.�xnT�������s�WVCv^�����*{`_Lg�uX��8n��F�v7]���@Wph5Iʆ/d57x��cQ��3����F!���o$p��]n���Sl�.�sl�����E�HR��,zu�Sk���=��)�A��:��;ǣ��{��%����@ b�(|6�A�y���|T̮�z��B�`��ġ����P��S��(�+�X�N��%e���dj+~��C N�,�/������>���$(۱�T�w�0<,�Z�L�.���匄_ �0*N�e���v5dh��u�zv�A��r���!^J�f����F#�\�V�8�>��5r�/z{,rz�\�
������ŝn�`J6KZ[5+VG'�R��*�YQ@�;�䃤�y�)Z�I&\⵨Q�P���廕L���K��u�l�N!�;��O����� N]��-yH�M��Ƴ�T�2�������Y��y���yS��?�g�=7�Bk�ݥ<�����Z��2ɓg2BC��+�� ��%������wPy|h�Yaڸ�]�G#�_��7�Sǰ��a������$�Bj�������}��4)��4j�A�c�xz�!������sB�`̭�#�U��ŝ���'G��EM"����N|�Ɋ��=\�R�*�?_��p��<d	����&���`Q`��g��'sX�>^����q�Bt.v��+��#������ 1P}�4X���'�U[�k?�G^G�^�S�𥺥�8t[�+~i@������4���c�iV��JBu�e��R|�P, ����%O���^7c�V�����D|S`5spظ��w �l��0��t�l�%9���=ZwjJp�K�T!J��Au�s�4�<�њ]S�#�x#�M�<��ua,k�CQ2��K��̑��2nj�>��޵e�����P���Q�?߳v�_s��L�T�^ȩ�0�ñ�Ӥ{���#���"3������|�Ϭ�*�x,N*���؊�� d+ֲ��~�t�9d��Q�@]�|�s���>2\KfD�4q7*���kI�����G�B�GUuϮ��N���6u�S���(���q';I�L������S�����D�0xN1�+wS{���^c�����ou�3��i����Mu�dq�Օ#�8�W����#�x���o%��[M�H�0���D��|xX� Ld&����]���O�nM9�fO邰���{� 祐{������P��>b���U'�o-_yUo��]J�z)��-��#R4��0%#= ��B���R�4lU�:���!c��wY��
 )sE�gy �u{��}i�H��~5�N�
�6�/$�z]#��Bxւw�Wm�2����<j�g���
��2*S�M�x�����ߘ�:Ц���S���~�[74P>(�� 9}�Q|H.j*FTN�����g2��F�T���9�rs@��!R��?�E����V:�\CpT��*�oя�%�&��f�����|�f���e�+"`�����s�5�Z-%1<������gZ߼�.�O��d���$�K��j�w���j���v�]L�o�F�����J��$��f�c3�j�,R4	x"�t�x;T^2$��R�o�������o��h�"�5�X�������/J�2WNU@@<�U�N��A*�F�k[)Oƪ�}��]v����"�'�6�Z���Bx
���߭{VS�1��^(Ú�''K	Ӊ	�����y��ӈ�.�^n&՗TÓ�,�xj~콵�(��x�jl��#�T���l�Zи�'���:���M/��"�w�c��!����|g���]�%�H ��%�謯\b�40��+�U�P �������8lVz�r�L���9>:���8�@&b*�6_��⢥�,��g;��k&�n~�g���l��[=oS1�P�,N��i|>�P�:*����g�~�<E���l���g�7�n�N�Z��M��[��{�
���'(M�^�7∾��j�_��L��~J�kk� F$�\�1�+=@�Ѐ*��[��q�����eg�v���c�*��*Wz������з���*���7��z��e[	��G�Y������Lmd��O�^�{���[�
pu�9�!S�o��Ӽ>Ǘg��E>z��c"<����4�V�������O�Ԯ �l� ��<��F>�P��4�c(f"�wT��N\�Kk׼���I�G)���r���n�D;.���ρיL�/�z֓)d�����y�#��I��<�w��o�/�Ǧdq���8�����Ea��z �)���yU����G�,"؎}�h�\<�0��F���Y3��Q��E^X{{UrsE�����j��xO
q]a�Hw()y'��k3�	���3���~�vu��<�\��7z��nίB�y�]}�f�q(6�<|��󌫹�ë)����WӎVl���C��8��wz83]��wW��'O� ڞJ��P���X�WGKhX�mNJQcֈc�{爌��ޘ�u��Yۖ��a�	x�
�vv�t�rR`���\(H�`�2�ro$#PYv��"^�&R�]Pd ,��)�X��{�a��LEë5wC�i3-N��PT�
�#�J��_�?�4;��a�Z�����^�bJ�o�o^~-I���ęD��CG}��	���T�l/�	�h'0O��9$홚�3�}��JB�>��n�Ry� �bO-զ�<�z^�i4\M�c���`�3%%aL��Qxj�˘kQ �ǔ��˘��LVr��m�m���o����!P��e�6� �1ߛ�M��lF�%�8�d�������1�Z��g�o���	Y̔���n@�栾UTZ��d0�����8������3�5�+���u�޾��L��}~|�������uO�,�������2/�O.srs��W���9��b�9)4�ד�-�]�!M�����ߺ� t�R�n՟�b�6����#'�[6f�%<�"���7����(�2�!�Eo��7v�}A[�N�P�:��N�3�'�T�a����L��V�/�,5w0�9Ϸp�:,Qn�M#J��N��qЪ#�B�������A��,L ��h)�{�,��}ۋg�T�(91T�I���wy�$�(_����Nc�r]��#LB�勖�(�����iW�?f����?�!�h��Av��~������F�G���	<�����u�b~`Q��x��4�I���R���$
�S�
쉕����4
\��~�����kzǎ ���6���T���*��S�G�����d��Q��|I�d�U]{%�;��\9y�A��F�A���c?g���������5o7����,I��f��s�Gֻ|a(�m��������[XQ�*�Ax�����\dVF�p�>���E���ǈ�c��'��r��6[��PJ�@eE�6��!m5��XÇz� IE��/Q^�g�~(��>����^���XUBK�!Y*p`@��4c�N.c56�%W���1� w����7,`��Z�\�28��>����e�B ��@5����w�T���(�Gq?#\S�3�or2b�BT��1�+ƭÙ"� H����Y��j�pq;k���-�u�aHJ6���q��?۠�=�nە�;=;�����p�E"��������ۊ�zu���s%���6U~���+ȕ4�5�4�@R��:�8m�3;����'�,J�g���ЃÒF���g�A��+"��tDQ�ֶ�3�rջ�����_��q0ԏ��_XSM��T�;�zٵ��e��1)�yo:��%���L����7�"��jy=6��RDnl?��8�U��p��
�(G��z3�� ���em���}���υo�b��
����$�Q�cb[Uc� GD$��ɏhh��IF�]�3p(Py��<	o��s��\*�K�����zg86����z�l��3��#X����ir&2Z$n�vVW�w�b{���ِ��aW*$Я!I�Kg�6�H�ȷ����������W��o�W����#���~��[�󦚦[㖚r҆�"]��՜g�a�p���Le/��T��Z�	�F֯�/�1��% �@/z�
gl�dqA.f\w	d��ɕ'�O70J�Swsc^@4�l6�Aw.��?���P�M�õx�ҕЦ ��K�d���y>@��e��j���g;Z5:,P/t	�Զ�[�;��2H�M-�V2)>��XI���5N��k�&�XB�N����G�}j��Zz��Uᘲ��x�ݖ�Z��f��Sei�ș7�+N�L6h�?�#g��"�����cI�s�5��u(�V�=Hr�e���>��B�P/1-�T�� �Wܳ-��5�c�ku�9�m��.8�U1�0��;S"��-�z��qG��;y+*�WV���K�D�4�s9Z�i�s�s��ǀMH_'ӦH~����:k�>�^��j���/ iU�?�/�H�
|6uLVt�{��}��>��)-A=o8D�L�n�k���D�>��`�ay>-))u��C�p�D$���
h���?@:�D����P{�c���x"����.7e��8��0�o�"�n2h#�ҩ;�%_bӣ��G�Y4�
6�s��Te��.f�kN����?��Q Y��쭰!%�������|x�&�;v�_�4ߛ��6���2�4e��;�xȰ�����6;�"9�ڔ�1��Qwxf�u��!���'^�a��h������h��;s�0�.۽�ܯ�b�Gt3�,9;�Ə	�c��%'8���cT�vG��a��z���w��/)��ɞ�0��S #�>'ꀓ�=�����Q��OrkYj\D�n�O��Y �aԢ?�UY<�� ڰ���':�5썽����wG�D�İ���Y��G��u!��Ɏ���~�@
i!6���*�(����&3$�j%~�߼lo,�7�6���q'&��m#�Zw�P��4ņ�ꋈ������Ɗ���� ��)�y�)�?��BQ#�9�/e����j��S��$I���-q�%�Q�I�� 8�'�u��	h���da���Q��I����E�37��'%�����Ǽŷl��G��vA+�������z�]{ȧ�7J�U�mmzYW�,����D�2��kuG?Q&�J�oz ���מ����u9p�&v62̕&_�	p¼�kP$�|�(*Uc)G�*f
$5C�O���W�ɫ�3��S>eA�Mҁ��n��.Bt)�m��;]?�^��ݖ�-��m8����M@K"I?>�Ms�ۇ�?c���X]9_�B��S壊�V1�m�U��!$A���2n�o����E�W���u�F��P����\m��F/�d�)�K]�����_.�"1e��5�l��/��E���Pk�V� �o9�8��ԩ�ߗ9������UE���k��ç@�&���6�����q�8�^z(���[�y	S>�vD�h�V��ԛ��_�SN�KKk9n��^���d	H����%���.T�(�0k���ʵ�Fl�i�Bw�"V�Ł���Q����5/
8Dfw�gAG;)��7E�ў��ѫ�������)���;�tk?���s��g�
w�L ��E��#�	�/-�a�@�o�i��No8/*� �9-F s�z�\�-<�q�-H��t�����W�P�=R͢�]CZ�W�F�P]�<Z7�Q5lXwW�#�m)��@��P�uh �d��VP�/�<�rem�A���"�vY�1��[�H)�n�����O��j�@X�)�5�_��z�k�{�S4ʜ��I�͐5�H\׺O'��s넍'���0%���h��o'"�j��B~���)y�~�z�1$
���� �U3?*L7�-�.؁ް�`����F���`�OP���5�T) ;���y_�词�|�&�z �Ljt���*̮yo}�ú\D}]�q�cށUqT�$C?f�kn���V���R�U�M"�c��T%\�m���t<i@\N�}�uF�m�
��A�2E�!���B�ټ�Gy�rt�\�iQ�����գº`z$����?ޗ�\�+[��챓�gX���f}Y��Fw��T��rZ%����@���[d^ݭ�O����.e�rn�lf_7������]_�t� ����d�0��j��|��#C3����D(~Ǧ��Sy澿���]��
�&��ߐѠ�eE���������^�r����*c�B	ѭ��#Gl���W )K0[�;�ڱ�M���V���'���"�CRuu{�@v���ZP�RO�ˤ�j?Q�{�G��ph��!WfE"�y�5Vq'�	26{�Ƥ�ŧ��?A��)��d���Ji��8UG$Wi�2�0��e1��|�bn�U?i�B�/��N؜-Q�d�G(C�>�]�NZ/�&�_a2.�m1%+H����%ISx�y�����z�.!N|���at�Z�l���(�m�#�hD��(�WҌl@y�j�R[�]{R#F�U��,��	��i���ka�6C�G�ǫ�ԶRV�Ȃ������t�Lh
	{�q>��hI#VvӃȔ�5b�)&]�
8���������zwFr�O��V�aG��5����-�o�hۤ���ݱ�:.���)����,~}�����'�͋���@�rdT�
�B��E3o��,0��E���6xg�=U�jv
O���r)��y�_��V���������K���O�2|��fo����E�jy�z�E/�l��b�D����2���.i����Eˤe_�W��K%@5VΥx�%�m�O����M�Z�FO����o�j��tΗ��=Jt*�ŀ����u��-��8�����l�b��x�0=8���}��vb�2M<&Z���Kmp)K+�����@mxd�g���zWĭ����P�	�=�;Հ�O��hy��
M\N��8PMW�������ɦ�!�����e����0����mS�A���E8��(o[�W�S��b�P򸀬-Oϖ)���ߺ�Ui�ե���8�Vl`*h��ť���,��E64Q���♺�P��,��["&0�8&�u�"�b���AɣO}e�@��*ܹ)��{��X�K0w`��NH	eV7�˵���31�*�,A�����}c��@����������D��[{�b�m9��a�Y-�R��Aͽn|�[`��{[P� ��gŊ�^��n�_�>f�@��Ǽ����4�1�0���}����Y&�<�i���ɯw#w��p��O|-�*��G���޹<-��@��0��ψ=��Z�����94*'	G�f�,���գ�vցN�/��.��&��⠗�7<:��N��5�`f�)��k���7�E�K�q�5�|�\��W-�����|��q1�)X�r�?ͯ�P꺗	�f�]4+�K���	y+G��i�d�'>��݀M�3b�f_��Z�TQ�;r7���Tb]i���I�	��������&��� I�3>�2�.S���I��5+n�҉�6����!��2�S`�%�}�[&�#c�aE�pύ��߶o�u�i6
�vg��}	v���݅��]�>߾�ѻ��Y}x��^���X��D���&��W�K�vS����ɽ&�Z��X��#�9��N��'��ah�w>Gt�����Z��0�MLZ�ĭ� �&Pb�2�����`�t�?iб�X �J�r��'�pnlX�wF �����}o�3��72L�麇���	Ԍ!��βU>tM�X(n���/������
2>��k�u��1�����9}#D�����Sy3i��!L��@_+����Vi����V,�E���F�ĲK-���ʽ�z���,�C]5R�`�$f(JV���9��?gB�+���h��{AX}��>�^6)��ߏ���e�O=�2ф��bi��+�U_Ҿ���H�k�"�u�X�mPi�r�+�p�й�rɹ۝�J�=�gu�yT���MĆ��i��`V��j���y^7Z��_?t���<����[���a����\C�/��J�B��7���Z�|CΦ�៽c���Em�ץTb�ޠ�~:�V���3B@�{��!�b]����'F�g@ۊ��# �.b#b]���w����0g�aZ(yE���E�m�Q���FX�E�'����t3Q���]Oh��k�h������`��AE�A-��B�/��!k��k�Ǖ�%-v6f���13N��?�R�:�ȟ"���^�E��dh�g�N!�vğwwB����'YYAe��_Fy1����)G�
J-� �Ͼ����&�*aS., G!��D��ӠF����J�L�v�D��e�o9|�u6��0G\��f��h��R���MA��}�,Q�2b�%���4'ᮤ��Nx�Qخ<�m$0����:9\>�p<jb]�/p.<H�66h��?=7@\L/���|�^!�%*34��P�����F-#-@��~���G�������'������/�k��M���#��3`L"j��-R��B��fxb������FNZ3�����5����bc$��9��L!���v�6|�����7�2��u�[of.m_;a�VOt쉜�x�|ˑ�gUB�9p���3Z���|K�H�ta�ͨb�_U9�����ۧ��-��,�,�x��c��iej��lh��J��+�
�4�w������ ٛ�ϔ��Mʱ ��8�{��/��槨n�����X�G�亜`	eb��zlP�a�u���P3�HB�H�$��<���\��M�9�6R�Pj;>���zc���CPP��pj����&���rٍ�!���Z��L�v��4�H���`�� S��O!	�� 2n҄�������.��ʝ��m�r����"��Pn�Q!�L˰uw�\.�&�,��Eg<�B� ���K�����o�GU�[[��a�=��{����ʙ�P*�W���7b��R# ᑸ���UMX�N-7�:�K����$�X�x�s�NYW�@QXmfxZ����x�$3�q��}	�E�v�/�j}XB�u��J�~�g9�n��� ��ws�}zI��S
A(�b6��flR;k'�c�\�m����X�YQ��1Ϲ���[�z�7�Y���$\`gj��Y���`]�Q�Q�x�k'Ҹ�����$3��H�Y���P�q�9\�Ta�o6�{�������tP�Ss��8�z�C��n
���hn������V9��L˅4���Q�c6�|O����Y�f��@�O��g�� M4���K���s�)��N��r�n���!�W�h�l&�}Fe|9�9	�����3Ec@"��Wl/n�U�->��	e�ړB:��!��dL�n๯Vsid��{,?�{��
a$7y�3l�M4Ju��$H�)��g0ǭ�%jK,9�I-�94EՍ�:q|�WhH�[��.�v;:v�B��n7�h��̊'���9�C�.� ���\R[+9�5 a�ض�����x��B�d�f�����]��G�ǥ���.��A��r��Uh_�h�hA�����O��3�qȠ������|�C�����+z�p�V̻z{ǐg��-T��ޛr�= Y�S	���*��&�m�tg7C�m'�)Wp8�����ϕ'QSu�H�"7����߮�����<Zs x�����>�����n�"�,~���G��[ɿ3hj"V}�$k��9+���}�X�ۆ�XO��V����y��N�E����|��\�R��۾ir�B����d�n md޵$�';���,����yw��3�&�$����k^�Q$���Q����Rjxx����	D`���^Yal��BR�q��n��R-e�Q�-�������_,����p�Be�ἷˈA(���\�p�F�Գ|��dɄC�q�W2�'�W[8A<�נ���E��G9������U,]�(R!��{ժF�a���x�+���[frG�kޕ�}���jF�)Hv��(�P�c�0:����լ� ؚh�����4�Ϫ'�J�f4��P�dB��n�t�8�e����;���sL�����K�Ө�F�O���,�����95t�⊣+Y�������I���0�6do��~NǱ
�D��U�OKu�"����ȴuxJa�:�<�,�G�J���%Ix�j��m��\Z6�i�k5?����i[u;�Bu)T�Fׅ�Z1������yCW�b�V�%��b���3��z�w8�b&���<�ۜzK&���z;��;���f Dӏ�q��7�	H������Ψv-炊5X�)�1��,�G�}�Ni�=�^|kP��x>�0ߩg�ػ���T�杂�"\��e�0%���	^��٧��X���	�����ܦV�6ﻠ]!o)q�,&�w�c0�;ue�˻1=?��I)�p��	��H�>�\��Q���O�ޟ��`���`�8�<I�̖I
��y������1�\7�׃'%
��⸕���\~�n�t�ev}W�cndb�,/���*$W��� TO5��P��a0���H����6���P�J��m�D�{��Iu��N�ai�0����S,�cr�`l�
9���;�I�}��Ő���@��Ѡ:1J���	��ah
�*�i�ܵ�i��vS䡖�b�5�Z;�*,�,%���U�h��(<i�m���H����78���2�jP�������#ø��SPMhV����O:U�|ض�|JK�h�j�&��vi�㌊(���<�6v����oXH>��`�t3?2���>(Ls��@�_*	i�^�!��u_�-�CfGe+*Gnn�!¾�=��^��ňW<�X��~��ّ�B�,x�1�@?�����TC�"x�J�r���Y�s��C��^���a��qք�E��Հ�V�wԂе��óW��������ȭ^[=���}i�����èǎE��\2���Uv��b-*�`�,
L�����Wb�*�g�\��qI�|s�T?����p��UU��>j�F.{5B�}� pi��D�ʄ7/�^�eԫ#��I���"f��z�c%.tO������kP�q���\�VeD�/���m��X�����3*�x�b�	aa�y+mxl�qK|�'�	|�Zo��_"5g~Y�,W�Y%bd\���M�q8�4����RfH+]�8˱���k�	@2���y�<~Tꋎ�� ��Q��כP��s�!@�[�[��Q��F�&��=�v�y�
�z�JR�nvC�MO3��>�f �E:�:�V-����������`����(��D���k�?~�5h�/��ج Q���	���%~H���uo8۳\������<�����<�r���H�L{�n��Y�$S�+P�$�7#����`�\���vj�^�Xj�z��0uq�F~�����*�l�Nlh��
��;AxR�ΜH7@�%�9<�HT9�b�)Z�"�r��.��]='���y����0����Ҙ��v���{5�]���f��)����j5�`�����I�������� ��A,Y-��4�|��P�1��%e����V���S@c&aqnar�A�D��=�vj𙀉1�|<�
�"�m~xnx���ݯ�~[ ���2�Z��V@'�^�ݵǖ� _frА�k��.�����^&��c�f.��EA�ㅁ�U�!���Jx}Ǵ��=��l1�����T���я�}�Q�Q�)x�2t�M:���,���\�@��W��*�<�*��䴌��-NS�D�h�6���.l�Us9��S���,�.�@��e��hC�+���F��3L%-V	q��/�fk��A���x�?�T��|7�#�� 0�V�Mo��DM�
����"7͏q�\���~6B��JJ���i
�����r�8 ��H�>Hvc�.)^�\��\�^S�D�CAR'��DS �/��mL p�t�S��эC�~i����� 
�AvD���F*��6�& �+�.rWX�#Hl=�7CYA)�>� �mz��&��\������o���Q�/���p�Z_%_U��ވ��e&Pk����w��q��`Y��6e��rI�����������d$*����뒾��UV,5Ή������V#�����J�ď�	D���IĈ�&li���P��Zc��2��jJ�3n�	͈��W��~���+�����4����RfC��2*��z���Y)a���r���X`3vЪ�q�B��3{ѩ���a��N���P�n�n������?�W5j���^ٕ'C�A����=�'����2���>��#�&�S�zd��;�"��O5b��֟�>��@q){����	�@5�[���ep�x=<����3���]��K������ιsTY�N=�^ӻ���z���;��%Z6�!j�S����f�L�]})w5�����ah�@��[���ߋ0��vJL�2:��FK�D̣s�M�����`�j��cǍ�=�G �2f��X1��t0��/iNi[ބq��<_p��H�'y�x\�O�L>?`�yG�/L?,/��#�D��N��*�q��J�l/�E��5���|?��zɨ��:�&��?TO�a��|.�4�]�
�6��2����Wن[��9c2��6��)� �{/�a�r��A){�|+FPID-h����Q�j�b��]�C|la�|���6�Q�oz�|��~ ���v�:Rʑ���W�$d�&w��\�?����A�h��'١�on	VWX�~�g���}�����L����WV[�9���9COB\�X&���޴���%	H�#�h��hv�ô���?[CmL��d 
H}���g�Sa|�F���9 3W6�����'��!$c��� g�Q �/�_����Y��`H��66z�B��ؠ��|	�.b�qh:��j� �jA,�am�L���DO�-}Vտ��z������\]��������t�=�8�Y��"E�����j��Ƚ;�}��k��2*7Iۿ��|�2B*^�U���6Ʋ���<�Ag�ض,n�W�X��4nJ�[��?E�O���0��rT|��M���LAp��.Z�ҍ�����j�5����,R.Hچ���5�c�F��j*�݂N���.���#��R�f�k�����շ,��:�q�Zv�m{��A��5]���*��Q��ȵ�.��;(������i#E��?��C~z�0%�������ϩu�i4�r@�L�u �k�t�:Q��ì���Y/"�Z�<�� ���"�H�W�*������'��UKR�0]�u
;��"���!��X�Ȧ-y�*��e�����D��꯮8���.����:�׫T�F�|T��Kc��-�x",J)��N ���f1�U]����6�'Ԩ=�f�J^q��J���;kyDX?�uETEQ+t�,��� �G1�p���5����bc�A޸�,��
.˵%t4VSФ��e�M�qE�5���i����Y����q��k��;J��.�gU\�$'<�G��T�3���Ւڴ��vW�!���`7�s�xrl��������I���������)$��L�2�iv�aO��!A�q����i���n8���â��ң�>ya�LGwa%Ҿ�	��1_��^@�X%=�~M^�����3�I�+U��5v,��Nɯ�'��!ЀK�qDr�E��W����^4R��M�;r[e�:G)�HҁW7 ����h"�����!zN�����[��rY���+�n����\��?���yyt"]q�>U&e��29x�|�� ?��נ�L������D� ��@��(�=�B9�j6U�P�M���T�5ˠ�T���w�O�t�Q�Q�����wm1��T�-��3�W��f]wT�a�r�l�_U;:Q=�8ؒ��-0EW��=����$���B-^��_�RV�X�K���'�ׇ�&6�he�����j�|��s�r|�M��΀�^��F��[_�n���uy��	ԃM���X�w,ʏ�֏=G_,�bd�5��u�ŏ�:��0�����g�e�&�o�=ˁ��D���q�%�+[:U*G��D6�l����,�{�˛و-��cw�IE�'|w��������_���;��U�_ O���*~b�%����<��H ���b<ͅǁ|κ!���5���6�Z���%K"�|@���ס �XT)CaPn�T�Zem�O�V�$�YՎ�=Me���Y����&��0M�"==���2�!]�=������`+,��D�ݮ0"�T�����	)K�si�Vu�-����k�C{�=��{���ʸ�Y���`X�-Y�Qs��:��q�^Y}#|����Є7�w�i��G��U��+����_�OtW�{�TvT�S�&du&�Xp�:O΋�T%*&0,��*�ze�/���d\욍*X���M��[��[���PY�P������DW>Q��,L��_���pp�h��� u��Iǵ�i��^$��.���UI�����-��l!���ybI����T9��]��������T��3�)"#�ςY�-j`����,΍:u�IM��[�@!
��ۏ�Ёv���ȹ��W��=C��6��a7H,��p�tG�m��0:}kޒ>��n�O��ǤA	�W%݂ٞAU�m8�v7��JBk�C�r�o3�2��^Q��?#��>�h��0g�A�RK�)�LW�&oF�9�t��q^���^�"�U)�{`Y<SZ}��L(T��ph;�����=�K"�R��F�D�;ܮ��A���Veф(��kQ���_� ����U�&W��P!��eWMQ��O�On��o���+�<�|�S�j���¹F�q4���	��H�������Y�h�1?#���
�k��u�3�A�'g�q��l=�ᆔy� o1!8� ���t�a{������'�R�t�HR��F����ӸJ}%:�υ.�j�������8�vԶ��B	9�e����4���
In+��tq��k�U�?��x4�1-F������+@��6V�'�)�|j�ݼ׵���6����p6�lqٹ
{ �G����+U�[�]���:�ퟏ�!%_�W���!Z6f��|?M��Fx K�g1��7?z�� ��Ē��4�Ht�R��͛Yn$��st�ֳ����u^R>���7SSNC����;�ֱ PW(�%��p��4�όT���(ǅ�� �_�*��_"���LD<j��3�a��ya5W��^<����B��.d3�WY�����R����(W_ש�i�(��j��<��M���ȍVމP�*�rC����X�Z�$3n�ū�f�g����Ksz+M�Ra\A�\�4�����&��	=�u_��I��"#l#GW��0ԕ=}�7��`X=}��Hv��B]�@�迼��K���.�N'��,a��5�Ds�������~I֖��b?�ˬ5w(W�W������-����뙴۵I<M�K����l'Î��͏���u�u�݆�~�i�����կcu9p?묩8Ll��{�:�VO��4��ĈP�N�x�,�!g�	\�W��q�As���:}8��-�P��斱B��8��ߴ���O7{�������xE�����h�����'hy�z;$m1����;��*Ilg��!3;s�]���n ���sB6���1Ll���Ց�"��	����H��c�Nd�q@?�g1`,a"�il�)�l��g"H�ۣ��� ��E�*���Mal�J�(M��/�~��ௐ1��'���z)H `�)U�!e���Y>}#���n-��4UΒ>!1v��*�N� \����uI�-�w��EBH�z�9�M�Z��Z��):	���1py�A����mWU��x�9�qV,��R��kB��&�ͭf��0�JFFjV�j H���,x��Qz��֌O�ݞr����h%]��Jx����]�����Ԝp��-$�-X��aW(
lc~E#H�2؋�ǿ�]�7��&��(4�*�8�����̼�����R�ka@�m�(�=)��@>�O��K�.���e�����Fq���e�P@����T������]���W�m�m�X �\5��'����]�6x�?		A4F���8B�ϵpH�C��TS���IW�+�0�@��T;��,����[f�J-e���EU7�^dټ�k"P��%ʍ�j�G����`
z΢��!mA�É[�f#�aP^]�~�	�a�|��l.:ua"5��0"�2�ݞ�c����*?���9�ˉ1�ā-ҋ��bi��?�q�86é� �{Ѹ/V�,���QD���O`�\��\5�4�B���x[�.��;q����-9 �X+!6���fk�6V�)38���6��lt�}"	��;��}�'צG���)x�7En|ȳ߶���5m�*�	N�gNz��|�;;~(i�Y�jX��}�b�=���4��1+��v8,y.DG����qU�7$q �u�����ô��/W�u}o.�6�k?������9��AW�!�R]\��TC�aoV^�-}�h�gRdp�X�((g��g�zL
�,Y��v�0�d�_3��u��#$�)�Z�%9�
-a����-�Lպ�d=p���-fNrx �R^��0��&�At��[���㰫O�|Qu����ţhsis��r`����S�����M^�툠>����,rwwx��>�>�B'{8j��8,'����df �o��.T���ju�D]o��J������s��(;o�a.��!�7�w,��A�"6a�\�T�C;��׳z��!���r��g����uF��Oø��/]�^%�_�G�94k!Qs+�o7�i�����\[�ƴ�QP��Y����h[�QK	�7��lF�,r�����-�Fs�=J,�T�j��&5���I.2�P��� �8?٫�.��[���4g?0'�O�[�_8��T�pV��%{(����δJ�KN��̽I�e���9��k���������h��C��f�R��|�ǫv��r��|''�(���B���t�;2~ ӄ�&�:Lt�tc�,a�<L�X ��o�f����>3M�́����`�kU���P�h��T�\�+���Ň��𳏺���ҿ��Z(��K:���ؾ�G
+}f�����Ų'�����E���t�m�8	p��
�1�3`ա�lZ��Ǳʣ5��A�KDS\�%���-kIOܔNG���-������swYai�L3�n/�� tS8��8�_��B ���C���\k�T���].�J�'k�a'���/�7�˝�Yٗ�\�^�S'ކ���H�Y���uB-[\F�����(�m��q�u�Z�ul}���2g�j�������G>ڪT��_�k�*���7<��ѿ. �^`f�p��S�&�9P�3��P�G���GT��[Q�LB� �!$�`�v
g&���Ln���F-j&��x�-� ����L��ܾ�xXQf����]	����yq�ܸ��{�n�^k߃�aZJf�9��C�YTB��ci��^�ja@���,_Z}O��P5\�C��;���h�Y�����L
���U�N<���N�yP�uMyi�O(�8��XF�Wz& �dt��j:�����ހ�)�D4�|F���wF~g�j�ۧ���7%��e�yHG�?���t��I�a;�ɪR�!m�ϕ�x3�&���|a�'��R8\�_\��l�Wr�1A?�C�(QRnzר{��Wp�d-x D9q
��k�[��Z}��re○. )�E�E�?w,޷fH{46��؛�==�sNZ2�52�5A���v��C
NU�T.��{sf��'"6D���)f�պ�s�S�38n��K��҄ͻO�G�H:��+����
å��g��]����L���Ů|~�ZƎ)���a��ф��u����d#��gL<������}��j��ӈ\��xD$}�	�v�{݀����(8�I������#�nEq�WeҌj���f�|#߻���3��h�g`0TI]�G1��^?��1�y��J�L�%����ä����d"]:�N &/2i��C��`ys�V ,����^,[�?�b�	�vd�A8�7�N�I����y_�̑Σ�Q��:�E�d��c�/���hoMzgf+�Ř__�qAT]k��	SݻU s���\6@�3�N~`�ʠ|y��Y`7@�av.��	�����Ñbqӷ\ʙ�.�$���|�v]�+���i���d���V�?�&CZ�U�p�c>�ّ��N]d6&� !�&	7�3+_���~Da��(n��f02\�DFSߢa~��^7��C����R=�[!K^��r{�EŖeg���K�+��\��&�$qU�2�!x�wvJ(�qb$n�	�Q`YE�K��$���l8v��$Nn����X忙0��:+�.Ji۸+w�l:U
�*[
����P�mgH0�,(om�d�YIo�A׮� �F�a�:T�R{�>��ag��r����e9�|�_5�f?�%\�x6	-p��L��hg��؋�2ؾEW�WT�T�����7ii� b[��[�s3�w�C:��RF��9��ar,�Z��ѤG��h�־Lf��w�Y���[��0B)ӫ�h��Դ���7����'�T@��$9g�%j1^��8�P+6d��{�N<'-'t+b��0��*Ш�eF<�R��Ul��!U����A1��Z#��Ú��͒����gfc�U�䕱VuU1	Oz��@)���fq���7�i�$qg'��22}*��]92��?kA�J��_q��}�њ4T���'�ߎ�:VU���,��9��pݔʅ�AhI¡6x�"�| � )� !�k����:��֛p�aR���F���K�r�e~����D���mٶ-�ښd�{��d�WϺs�|�5"v64D٣qVW����b�p��a�b�⧍���f��$%]�=n������ �0j t�	[���̈́�-o7)�F��#�r�Ŏ�v�Q��� {zة�����w�DcKE�ͪ!D,́}a�2��n(�|F����=��.���צ���x�g�ڂ���]��H�(�����e��kX����������qZ�CS�l!�,�n�90���ϐ7u�e����8��^���͗�i���G7\ғb�t�O��ҙ��5��s;�-'}Ƌ2��g��Cŗv_�g���$l����G(3�Sqn6w?���w%��Af�z܈������_Ϙ�$����%ug��GN���毹��/�����`3>��٦����c�IZ�V�-:x�4�'I�2��i)��q����4B����{M0':�[9 �EV��c�;�s�P����պ7@Y&$�ՕB�j�,	�1|i/��"��9��ѥ�$�p}uRՉA��kO�����5����M
;��Q�B���.��˘�� ��lH�bc �75��8Ѷ�$7�Z���~�w/���R��2�d�P��vX�'��X�f�y�A�����n$V���O��ٜ�A��8|Y�*m�ae�ᙦ'��i����#	6	�5�{q���z��~�	�P\(�������]� 2�����<�~�������>�qdI�o��x5��5 ��x���<[�?D�$�C=�ϸ������_�A��8}裖|������;�sx;r�2���c���8�;~�/M~��5��%�u�N�H����璵[�$�HKʔ��=�-��D?US���A;���b�O��������W!�c�l�$�Z[q��c׬]�q�ٟД��Y4�'����g�Uo��S>L{����o��^cy�m����8����/��8EN�
bA罰zÿc!�C�D�����܀���U����N�Y�I;V�^у%'��Px� L��=�}�i2��#���E|{��p��RcQ0�G3��1[��&�N�@Ry��b�R���KZg� F��Fw\jR���ϒ����'[ܲ��,�LyNn���Y��d$A��Yߴ���>/TJ�@�� c�&c6Dl��%��@՚�5*���#��MMң:u�|�ZuV��)]��D?��q�i�M�~�!
Z$%�O��ّ$�35	�U]Ps�GyP$Q����& ��O�o��YH�%�����ݽ�i���K@5%Z#�ѳ?�6uô�K0�ɚ�B���g��N�~���L���e`�4�sr��wߪNf�\?���3-� �H:����Փ���\&�9n�G#�Zuk9�M}@UЅ��YIcuO�\�1��j�k�9�FD~����Y=5���cz��5�F�j:��%����y��V�jl�ow�@z��O�������yIɹ�r�7<���7+�S;!�询��z�1�����8����-���T������\�m��4%4�:C�\�ד[�D�eU�l�F��:�̸�dj3#ŧ�1[u ��,ۍ���"��@0O�������K�G-\�j��VF<��f�w%���l��U6Ϲ�̩`�uw2̃X���!�x��N�iS�P�LE�Q���^.�#������x�Ѡ�GS3�D�<Iv��\����ա�5��S7��B�ǀ�?��JIm�߀��f�K_qW�:�T!��u"��^DVp	�p�f�W�vV+t#�?���f�_��)Cu��2ثwΆm6�اl,�.P����Y|��d60���$3&5$�y0���U�{VlP��&t�Ǻ���le�PG�����:�$F�(4�S�.��(�݇4#m�.��M���  �k�,��+�d	tnY�9�3"�ėP�q��>W�ʎzi+�]��V�ߥ�e�Js�G��4l��#�?/�n[]��8�H��j|r�kF��,�މ�R�o��X����fDH��t�o����Y@/����w�po_wW�Ȑ~�נą"ې�K�=�qS��k���%,�P�@n)?.5�Y�Ŷ�q���F��
-ٗ� ����7)m�1e�+oZD��:7�����9O�����?u)�v�Ҫ���7��_�y�Q�g����"*���v! tM�?l����';���21 ;-���� ���<CQ'_ܷ�{_	��$���^�7�R�0~�5= h�r�YՑPh���!~%�WKaQ�t�Z��1�Ć�ʍ�^��T</%غ�n\�����w�f��&�lޞ�(��q���� �&�f�� bPX*I� gA_ڨ�H�S	E����Ig^/�Ѣ,&�助 }$,�v�����=΀1�/P�3���^�=�+�Ƴ�5��wș�y�z
��$*Ogs�h�F�����[
z�)�uj{��0O�T��si�C���|6��ru�D$���[��鄙eB�S��:e�S&DH,� ��'ucr��v;r��a-��<w:2j1�!]y�%Yq�Ue<��ح�����:�$�6���$�!H���|Lj�NR������}���eH�
�koZv�j�,�Y.��'"|�m$��z�R���i��.�4�&^��$m��V���6c�Ƨ{M�^�OLsoA�vyqo 옑Sc�]�;�=�o;����]�Y�	8�]Ȇ[�iV$�n�ꧨ��
Z`޼Й�uWF���9�:�f��nT�s���5�;KE��)c�\x=�5��b��V��~;FQ���u.��4Ⱥ��6�:�e�Cq\��ʩ��C*�'���i<�n@ab0Y�������{�X"�]��c�X�|�*���p��h���m_��(�E�#�q˵O}�-(Y���M�a��D�cb93��$;6��{T���Lt��U�b�&�Q)�"� ���0��5�����h�Q��L-&��!@9�j6���dC͟�H&�5�f+�ˡ��>5�r9��<�+�a�Y38n��[��-� �0��&{����O#�����a�[p�v^���Z����YX'���9�\�m�R���� k.������MCSlrW��|q�7�� E��Eh��%	B������#S���tX�/����9�U���S�2
Ɗi�5F6��ใ۶�N�l���R=����Y�� �����ξ�vtZ$u��)X�	��G�D^h#�_lC�I���xт���!�zD:Dz,P�!U	[G��6��)��x�1�&�_�8z�4�-v�1�� r��mH��EH�Eɽ�͸>�{���(�LnwL��N��g ��Sc���~���Lh�{>�Z2ƶg
�˷�t����e���c�A��wN�x��w��I��̜��o8�t�����룈�4y��C9�h,<G*}�i
�,��c[ß�_[�`�7��~`�,ȫ\���g�A�ĭڂB��}����{�T������!%5n�I�q�x��@r���RAv͋$MLg�k�s��&�D���nͱ}��rAvW�d���ٛ5�}�X�DE�u
Տ�#�MS����M]��"�S�����3���!���'��=�!�LaW����9%�˷.8���)�i�L/ˏ�b��L�%��Saq�y��&��{]Tܶ��-U](G�$�K=��74��ek�a�)S��`�*��(�pk[hz�����Ǜ��H8f�J�-��Y�{<�z����`�B�Q��!A��]�(wYFD*�ro��jD���e�̀:Q�^$�Y8��;;uEo��;xty�tO����ӄ��i>3aq�����Ah��6~�𖺀��t�<Ņ�~��$��X��
�GA�Ѭq&��F/�N/a�T+��U�eI�����ޢ=5֔�Y~3�K��a�	�ҧ�d bR���Gfvp-����q���M�ğ��	�P�{"��:�Q�b+���� ^��]~���Mfa�dSr��ɉy�o�qa5S�,�>��̀L�2=�?%_�ÁL�>�b#�a� \%�_��������������}+a9z��HD�P@�gx ��]��3� y��E�������2�U9�+��X{��HZ��ޒ���Ͱ�����j�I�ȁ��wu�xA�'��Hx���J�x�� Ӧ^<9o��{$Y��%�$�{gN��U�|Ԯ��NPw�H��b���d?�N�ɧ=,�`�� N.M��7&u_Å������DP�ݵ����k�K�8�[?S��'^�ݖ�A��?D���OI�˰ @b[�e��SzS{�J���L��"p�t�D��M�!#����C�Z�o�p�s�B$9F�F�ӆ|M{9���3'��S�N���Өو���y� aYE�ͬa�{���)n���;c�NI1�c�7Ѱ��W
��E�H��o���� �Be��õY&6
	�1�(88@����Pa�bm@�W�Kt�ΔkXt��vv�r���(+2�:��	�=�;G��fB�w�?[b�_��� (�3 '�[ݎx���v]�Ѕ���~�T9�����4�y�cu��J�y����%�9��ˡ&3�^t ��l���t}b�ў���ʿF�oyRG�c��X����J����֨m4S0�.yu�A�X�Zs^��\��#xBxT2]�pєG�c-% �6�%HJ��G��S$�F���F�fK��SǑ�ȿf�P;�m{F��`I(�a�
Ꭓ��MR1�lAq�o2�$�Ϭ�O���4��
��������^�2����a�L�Tm8bIq���O�bc4uWKs9�M�6_�o4��^��ê#���Ʉ�P��4�Ԟ^ز4���1s��ŃF(o�����;����o��a�Ҭ+z��܆c�Q*�c}����WߢԌr���bSvPbu�����z�0�%�s�?�b�O�T����M=u;~�����	���!�3���6�^g���Zo&�a�3�&��Ц�r���K�wi$�~~�5?W� �zA��y!���ԗP�[�Ց� ���/I�.��J����ڃ�����Lh^È��Ӕ�����{ؠ�Ć��cz�S(��^��PO]��tK�D�$�/����r}ԓH+�����ݹJ��SJu���P%�Ҹd�fɾ����v��f�9ϕ�hz���~���T�-�1�B��u�吁����n�i�vI]��r[�4�=�ъv�*��,?���]n�G�|3tފД2����]a��eE� ���]�8>X��t�r�+�����1a�m��u�\��R�1Yt�7x���L �����f�q���g�rP��ϴ�p��xt�Dg�ì6J�J���u��4�%���?Q�9�i*G��Ju���da4{���˔�J��T�.X=���H��*G؀~+&\�Q��,Ǖ�� �wR�9�6ѥG�4��<���%Ɏ�>rW��Y��	y;��y�O����Ė�
@+h����)e��{�閇=:��}�ڰFaEO�탠h���= 
�*�V3��G�˷/*P�9���|�'�e�������~���d���h�s�#xGk�������������}�`9S�	�5�����}��~��3�6����wƣV��.٥��I���4z#�:���	���K'^��v��B��#�XD�.٢	(� ��=��Lו3��p7��u���dw���XhJ<5R� ���y���ɤ\�{~y�B��n91n8�!���2����6M���SD4~{�Sv���e��t��t�a\9�N�����I�G �|�\��U��{����@f�f��%03����T���G��������x��ۯ��Ns|!�RTF�۰d�|2��Y��@r`݇��Cڡ:A�2ի��M[@J�_~6jd�'P?N�(qJ<���Ä^�5�L��� ��1�'�-�ҟ;��j�5~0v�0��љb�š|�؄��O�l�� ����į����K�H�Ud��2h���t�Q��>��ge+��¤��%�ډ�^��u,��3���_�:���i�4E�w5��}�Le^9�tʚ�	��.�ɨmi���&=eY�N�#�j��6��C�tE'���&�Y��P2���T�
�5����tM]��g�$ht��]��6�Q&�[4�`����N\�����
p<�籖�/ C���ٵw��FpV,������~?x{p�C�p�Ԣ:�;�,���AN���/|�)�ơf{_�Ml�{�x�;�. a��F oy�-*7\zQ:m۵?�^��
X�y?(��e����J7i�k��"�1��� ���=T�t�~�2vA���s��>��ħ欥 �&����7��� q��^J��>�ކ�!LNSOF	~8�Qez�O~_ibPjH�(�8�Y�A-��w�v4
TW�w�,nx�t0�0�6�����,�4ٽ�,!Ws��&V��n4�}?��P��/���F�Mc'��!7z�s�O���ON��L�eH�?Bڎ^G��o�[�uC� ���<��H�C�m���)ֽ��8=O�f����[8��ٷY+�s�(��AR>�#L��Oo�t�GZ~ɵã}
kX`ŗ�n���p�l�#���c���A��-!�ВN�����Ӛ
��������nX1�U���n���_K�#���ş��Ǆ4L�f�!ˀ}�(�{�J�qkC���l�Y����1?��)X���.�Â�Z�ڡ�Sa*1��N?�I�,�+���֟i=���Q�8����A.q������(���J�,�i�`8!�3ƻ#�=�f����.�̛��\�\� o��QK��e.��v��"v��j<]��,���hӁ��&�͂�W nq8L�s�a���26q�v��������4���21�ݟ��b[7�x����J�r�J�;�l�Y��0>F����= �S�ކ0��K]ɀ���P8�Ɍnd
f��A�~O��g�~`ZM7��b.[���b���cb�:����rQ`X����k��z�;�u��h/T�G���n��}�41�������bCL� od�� ށ>)&�D Ef�~�\'��?�k\wʝ�#Lb��b~ٿ�ᴅ��$�3Cm_x5�:n�S�"���?�+z�U%2	��&�ؽɚtR�=Fk�90�h1����*�pv7 J9@9@ی1<.�;�!�lʰaop��iS�`KP�uWl��� Ŷv'Y([K'���!�P����b?.��$@��bn,��&zE��Puyߊ���p�V`%kWo]M-v�f���U�����+�W8��v3(��������O�w�,�='}��*�D&�/m���ґ�ԩ�G2r���<����QNI����}Q���'j�b'K?:�~,&����e�OSڤ�Z$�
��]�eNǡ�	\���笭�>�����t?�{h�
���n�<-�0�����.}ޜ!�^H�������Ok�Ar�V�w����'|���-�����_	����2���_�z�PtO�k_��%8�����(#`q�PB�[�n$�h㗞힚@��m��gB����Z;��gp����w���׆2��/s>�S��r�}V��ɾRް���zy������:9N܁"��G=v�aV�Zq/����EDl�V褅`u	���=�^U�7[`=7�N�������-Լ�`ܗ*2Q������[�#"�W�v��*a�u�'�Cv��S#������P7J ���,_�mHOQ����kg��XhA����5(�A���ROMS	�Ѓ�鶼�Hc6��'���|��/�!�j�ȅ"��R��"/%��X���+z`EZM�@%x���(@c4�?��_s��<|m�HA�L�6���Ê����N����tG*-&��N��ȃ얂�۸g��D��`~��X3����s��nI�׃���;WV�]�	��;��B���P��^�BC�#��ؽ�f�49	R�j��͢����F�8�̈����V���*�D����mM��V~\�f��G��
�U:BA	?������:`�� 2�Fn�C9���@��	lȏK_�� V�����d��_���@RϪ��@�u�:Oc8'M�,�>|;<׫M���-�T�K�e�b�Ҷ��2�.�
t������qůK��h)���b���ݜ��ah (^�b���$C<�Z�$�8���v��P�br����l�*��h��CP���u�"WB��~p5��ͩR�+����K�u1��(t��c����ݖˉ�����=P1��1�u��smna�P5���ƺj5Q���ǧ�6�z������@����G ,/��2���p���7�כ�����Vڲ�`!��mC�?{p��z�3��29g��kU��;!����JW�O�b�J�jRo���0z6B�� *�<����9�do�����h�]�\y�0�}����w\���~��*�*W�	#c�t&�$�J��f1��u��#�ڧ&��;���ы�H���i��f��%�p����s�p�(|#�������z���2���V��d��<�5��+�ґF��q���ӄ�K�gF#rͱ�0� �5�	dU�S�F���Ԃ�ś�F�z��ʚ������%B/�����g�t�V>�Z�
�'��&y2M��G�d����ʀ,��$_E�qU�L\ZH�'y���n��>3��'����3e�6�ܢ)|eN�HQYev��I|�32���勅��m���P�����ꀊ9'�m��S�z�'u<�oq�k֑���h���l(DZ��x��+8E+����+��t�;��s�c*�
�>��MXѼ$,p�s�E��7y0ND$t 9l���FT}��e۽�
1��ת۾U���4)��A��Ō��e�G�Z*.J�8���Tm�r�O#���!�R-�tM�-$3�o�H�C�l�]��=�0���M�f��P0�j��Y�T�3J;�֣�P~7iQ-�T`�Q�!!\�J�f��=�@�C��̸�6)���ܪ�#���G��J=��a��}ް`>ث�����e��(�,Z�MD��9�I3�	J=7�-I\'��gD�c>}�_���a�n퀧��Lݹ#���s��_5\C�MM�L���M����D�]�z<s`'g��K�g}O�[ �'�+\��}�s�u��?)�W��L6�$y;(�u�`+B�^>�kv)/J�0)�=7���V���mc�bs�u׻bF�O=�[��D
n���OO�%�1*���7�́%�5V).��b�Xc$�M��{���'d��p.��	N�ǒ�oөT��B��������Ȅ���M�b�{8�j���Y����G��p���P+R��w��+S
 o=���2P��J�A-T��O�:� Y9������]�>��5�}D��_J��]��vE'����O��,3[��J�o3E����� R��b�ڇ&�ʱ��=M6��޷O8h��gtw%��fs���m��˺�~����;�����"@�{M����Kg/�2ۿ���� �ٵ�{ �D��-~#� �Z�k���tǷ�B�wlX<Ny�<����ޡiR�[�;)u�{������	��K���5����\��� q8N�+X���P��G߼�ĩ/U�r++�&ϘUC�g��
���ˬ*~	�g�����\�6AhY	��,�w��7�x��6����Qձ�4'k����4�h������u���!���'8?h�ʕ��F`�����v���3���WǷ�W)��=��kY�"��A���#s���,��}�>����
]<V0\��6��Z�V �(�®Ql��Px~L@6�H�h/��I��?m��N����8�Z�����̸�]�ڞ���练B��tlQ�A�8�i��J|�U�eTon�ӹ,!��[���
�#����/��ɰ'��\�W�����p�1f��J\,?"h{B����2�<q9����Ȉ�V�@��TDF�ߙ�Չ����q�������9�n��	��h=�͞_��!�M�p���|#aԻ��i���QI�7��3�d��73zGp^\�@�gBx��IC�P�G�)s)�_��R#:�Rb[��i͓���_�u��JK�:��v�Ҍ��R�E�P��d�1�''�H���~���Ipˊ؛u���qJ$��E6_5�@b�`h�{��Ԉ�Kj��?, ̰�����1?�o︀e��EFbA�mEv�Sg�Ҩ��-�R��8���9_S�uC��},�Y���W>����I���!�: !g�����P��hAX�j#Hr�\J֒�hH�&L{<��a�7Xq��);���!R�����e��?ڄZ�_{$���r������	��a�QGU"=��eX�޴�f�3��ſ5�0aWt~�Q`c}2o���-�2�i�!� 7�[G�&��-����C$<R�e]9N`)�11��V���n-��i�U����2|������� UJsg�qu���(X��U��?���$d�>�k�o��J2Vl�у�F�1�xc�k^=�f֓Pi����yGNas_=^�B��k(;A�Z��� ����}�Jd8	N8���Gm��4�@ܛLL�p-}��?���÷�9��Ҵ��v�Q�#+�$g&X$
ː��,���3�����aw½�N�7-'3/as}�V��H�c��� ��&����t�IӃB��Ե�Т�_��FXUu�-��c?��f��mpX�aPx��t��,;�Y�0���:�=�p����A��A-��uGl���/���x��ￖ4>�toOS4�*ޜ���+�鶊�E�c�X|�T��\� ��7D���Dy��|�|d�� ��6z�ﺩs�&���5��ϗzoM#���Pljy��+D���}��6���lϩ*��d_d
o�����^�3E�u:2[c�r0�JN͕q�D{?H�0��p�~�!)�M�G'��Rz3$"�G!����������奼�WaG�ͨ9Ջt�禾�<�y�ᯣ�b��x.���3cS�[��G1��W҉�&�� A�eߴB�?~�ttp�%��^��2ч� ���/�f��\ AX,�+�Ɵ�	��2�i ��R�ul��������$_��J�/��j'Z���8bF&�tv��֐5��|`z��}>8w��E;����c���3`�x�;�"IGr�|�� FՖ����<$�h|x��
�9A�򱨼�*3Ԟ�f-��2H8G�PG�����^'������ٔYIo�4\*���j�ȒXX6����w�s��q��Em�Y5�o�np�)_ݧ��`�����U��A�/��,^G3�����H�u��I7�q��s�+j٘�ٻ1�����;O�b�'�|4Yԛ'Ғ1+m|���!��/[>�x Y���A��סXW���W�O*��sGl�\誣�8�涏<!Qr�'�_e�ż?	�6z��xB`�#�)�	�%��'A
Tl�(J<J3/h��8r�������zx��O�]3��{D0Z߇���wZ7.��kw�c����#��?��O1�֎����V�c����;���X(p�_P��X��ʭ	7���}7���s�ʊ�0����2�љxf/����)����P�R<&�|�BUЊ�3�B�����0N�L~\MǨS����\W�Yc{��rו�}퇔I�0ƭ�p���dd�$�4C���Mxwn7vOą��$����� ꥼE�5I���O�S��9k=ʲ���(�55�J4��
��Ldi��-��1Ll��WG�"�s_���r���{��F�Wگg����ZN��*��i��Z_�ˢ��<̍�<v���ۼ	d�I��a��~���[J&��L��䢀ቫ1K��*������:�8=Y��aQ�ǰ�9�2G��ϥ��� �m_���L#S�	������ _�G_���(B����Y!Ɇ��̬!�p4�'�tT��D>���?�ϕa��ôByև���nOIϬ��l�ڙ�x��j�J⣥`6�F$Iޭ�=;O���څ@V(l��$�B�p��A��շ�:��2�m�f�!��
����b~ ޗ�nA�[NR��ПF��P�����wZ��F{�ⲹ������h�i�K5~r���T�v�.���<a$~��O�O*l�5\�}�Ђ�m
y��<]?��-���y��oo��?T�[��F{L]����"��(�����(�.]A�ó��{Q??�"  ǰ��V�. D� �r�$Vo1��'oX�9b��������a�%NV&�_PQ-?�.w�XZ�}�z���3���crD��nf0cm�"�H��@9ޢD�� �%!fKnL��f� KR�d<㪓� ����C���x7���8��1��"����Tz��|���<�,^#}�_�_��٤���._����"cO�t�C��|=�ޒ����O�N� �Z�<>N�y�?Ê�����u9���"��Z������"W�I�w~��I�֯+�*���x��_�O��/
��)�'��ma�P~��p? A��O�2�{DT���Wc�Ĺ)���`a�$�D��9}:�����'욍�[���}1�w�]|R{��Y��,]��Ԑ)V���aR$�H^]/�y�DA������.����(�<���p�f.VZ���:K���)CWI�Pr�|��5f���s3��_�9�x���Nщ�V�A�0�FV���=q��z�Rk/��<����B;��`j���1j����|ۢ>wo�D�^�r~\�2�r9Ui����7��n.�<��Kv���k\�����-�.R�2��/�h��j5�'W!h
6���M�?��B�����S���R/9���%��5V�k,��u#B"ul��rG֜���U��٣_p��?�s+C����@|����X�(�
)	F��9dFRӉp. s�+�7	EU�c>~9�#��.��D*sfu���2?y��p��~ϩf�
��c�5��~�	��da?���4&<��]���^^Q�|�[��G\8�2ڻ���m�� ���h�u�0D��|^.�u(���d�&4kZ�B����=�/ -��g�}��W�0<��c[��0�4�YՓ�W�>��ۛ#����QPܝ�t��4ڧ��}�#���7�ћd����}ڰ�������f���dR���x����ZN�T]T��n"��{On�w|h��h$�E���8�NŪ��|���,��Z&$��>iIP��p9~=�ŀ1���D'����\��Aۭ딭ܑ�^v�]q(sG�+������v��oJ
pXW"SVl%�����jW��8���E]��h��{�fAF�i��x]�9e�R�~�����k����4.lsT]�mDE��@r�+�Uh�xC�L�ք�L�8�L�y��R|JޥQ�oK���T`;�9�1<Zm��t���fdt"Qc�H��"�3���˃���g>��5ZrK�/l��ŷ���5*�dǡ��x֜���t�+�#��I�,w�i����:�l�bx�1�c�o.>���?�Ŧ�����phN���`�׶O�I�bO;���x��G�t�M]�4of����ҏ����6��X�pe�j���PK���nWru13%��%J��Z����L��.�a+3�6�&ב0*B_J��t�L2��b��n�j���lZ�v{<�)R3��ؤ�F;g�8�6.�X�_��텵EA�%&�(Xtye�lz���3�u����X��R� k%�V	M�˘�Y�'RlL��d%�Ѿ����rK�e8C�8�%�+��0�xꏗ�	�#�ܲ��w�\�)C{~�F�>K���f�&������Q�ll��/2{�<RP��|��ݧ,�?�L��t����=l���~+����,A��bp�X-�f=���X��̌�
ߒB!�@,-���T/U�Y�lPN2�����F��������� v筙�P�l����>$��O�2M5r�bQY�Sm[�'��ԝy��T�tٽ���	>2��,}�т�·���31s��.m|������e��Ϫ�|=�O6�:dV�%e����wI�M`@���$8,��}���ƍ�e���e����sMsab��cU0� v�1��`7�BbX���"�� ���6lp�#8.�nt��nܮ�U�p8��� �rR$��J�E���m"ة?=����,&�(٢N���C��T�Hw;�r�6/t�^�~�u������_)ͫ�§{�������T4S���!�72?x܉M���T�Mo"��|��!�$o�%�۶L���?Kv8�3�����hM��K=G~��.)��f�mL���M�ݠA�C`,c<���y��:����h>��4>�v[�)�3X��	�Wz�Ǫ����hT:*�>��YgU����L��������m��$ؗ���t:�gz���}9���U"��r�,�vu��H��A�bf}-	A��������x��\����4������b�[3��Ū$���-i%��"3
[�X�Nh�-�o�bv��	'���d6�I�:9:�!k��"Zzd���\��� ��=����F)w����hu���OÊ48S�t�I�[�3��4�.�v<���B�A�~���u��
�d1l�c��1H���N��5�~"Sr�j4o��ap�tG�w蛔(�"&��?�H܉�{I>7q"�jNQ���l�,�RPxgZ����/"��E����!ml�r�D����$f��kŰ!6�#�̡��ړ�M��1���^<J$��?�U{�b5ϲ��\F��O)���~í
����2f���x9���rӴ�fy�`C�'����Ϯq�|��]�on�3���o���բ�a�"�i��v��w��bqk����oq���&>�C=�呕�"�m�>�CL�b,������ؕ���9�yao�f�i��R��\XI���LX��z.�
o?��|��H�)m�����^	,)WI���~ͻ�O���ϫߏ�4������3=x0��4����o�"���ݩ�U�JF_�˵��:\: ��Yv�����x'}�Y���R���U�l�i?�aD0���\��'Y9RtNqk�`��]�**���+:���fT�J�"9;Ͱŗ��&M�`PRq�I!٪ߞ�ǀ�°�㰜i�ۖ�U�M>�f25�	���	�;GZJ�I��g��F^}mO��đ�˟g�N5����"/��-��&��:ͺ-Kz�;��v ��_�����\�Z�Qg$C�o8$�V�wBG�K��X�1��r0�GW�1:t��oT:��:=��)������5g�&%Z@ �n���FO��z1�o���N :�1�r� �X� R2�F����x�M��%�%))�������������o��j���⾮�\�x\f�V}�+o��p�s�G`��oEIP'��0m.�47�{�F:�����2#�=߫���ȅ�l��L��:��!]N�Q�F7�$P!c4�nF�0m`���ï�->%���F���bu�竃n�3S��Db�ξ��+c(� "i(F�/��S�@�fa�Hd���Y��2�FH�(���]��z���A0�&�Ueb+?J��:j���Z���g��u�K�JSK:���`�0L��Pi��{��������.�$��y}>N��{��u��`��F4��]��.�Z�b`2R��[�����``�I-^����ITʉ��hCj^�t�$ �F}��~��DM���j�ќ'\�H[���3]b��N;e/�n����Ҙ��1`zu�&6RRK����p��R�G�spO�Ô����Q<D*�U>YL���拞�Os�׀f�x�{<-n�Q�B�����\ė0B�Ȱ=[+8)wnIʍ9����J(���O� W��_-�L��g��j�ih��=�e-�v[�t�����^�0f��-}��T1���p�8Lˠ�b�I8q�)�������t�N�'�`c�J1x�J���>��$s����ޒ!�z�71º��F��_:!����2�@����R�.� k`Ӂ'-|�!�����A�38,�	lv~q�O.�I�	�C�-!�3g(��)�Kd`�M*op6�+����@28>(�å��Kei���1	��i��̺.�c	���M::fA$�|S�x?����Sc�bfr6���I������u��J�c�������)�+��0�V��T4 ��=-W��������.ľ�� ��O!�ә�F����tɟ�8OըB��6�+�D�tXiH�ѕ[��tk�:J�n�����rd�TL���Q��%�?������P~r]:�'.ۊ�ȅ�>�C!��U�yq�ef��t�t����y*�q�u�do���N��} �o(��bӰ�@&�(�sw�������$ixM1�E�ܖR'JY����Z����� �Jz�{u,dM���xSlC|�21u_Ѷ�N�Ӡ0IBzſ!̲� �;=���c�W� �.`�b����v��O:s�aqV����R���G�X�ږYwW���s� ��I�Gx���I�8�zl~i�p�0�U�!Ըui@��#�]�o�l�����-ṋr��>�#�eȚ��Tf�$>�������nğt�7���^7�f1g�]/i���O�v����i��s�l�S��7����	W�Ś>NO#w����S�̓g^ �m�����47��G�`�Q�V26��+O.�R1eA��@��t9� ��<1x��D�#'���4?er(̢]ۥ��v��ƉZW|�њ��x����7��[S��\#C� ?���5;`跎��c�Ol6L,��ai�����==�u�UZ�Dۉ�v�36?VW��U!�W?�.<ׂ�gr~)�����w�����;�ǹB6q���<�8�]D7̦8J����b�����9�2x�r����,۹3���J���bM?,mI׳m�gk55�\��M�������_�ű¦�E.�U lGz��(�ֶK�B����|��L�����p��p�<4��{
z-K(�s"ˉo�=2t8�P�7e�3	y/�C9	H�8 j����,��BhںU�����'���ߣ�:�yԣ��|С�N݉����+����\�^ �ϙ�j�|c���o��4`����q��{��FQ�U>�bߌk�����"��b̂����:?������Q���PY��t+��2|��4�f���f�YjK�&��	��N!"L��g� �(�K�jM8A��B��i� �-j�[_C�s�"x�{!���v��'�)�	5��1�'&V�W�]���#on��ܾ
�o,²�L��m��;Tl[]Oޕ�R�J\.Jcؕ�c����z>��_���:�'��3yj�o-����&3:z�;��ɽ�VB�(�X���L�R(g�KCy������7�UT����GxkH���Ɋ#��^oؚp^��#�7�a�������rD�TRH��;�o���Ɯ^�6�~�%[Q���U_"���?�q����@��,�� 4E[/����9S�ԭ�Ei��Fw��t�Ԭ�b��r?��L|��cAr&Z3�UJ`-Q��7Np�0׵.�@S�Z�q.ݝ&D�x��5�1�"���>�6��۾j��MՎ2���az���[�O��rh�]V�2)�b�y�� U��X8�*�j�w��	H����*\��s"��-G	�!"glG��q'����Kd�Z�[�B������:e^ȅ!�*\v�z���g���fۋ���W�S���6�#�(o��7���Z�?��v����4*�t�?B'�?����SGu$6 &��λ���s�kU�9A1ϟZ�:�;�6V��G��2��#�kn<�I�r|���D#p�k8���b����
m���}��t��Ͽe���;I6�A.��i��I��p�k*�!P�hv����V�hA\7����Lz5|^,g�7�.}��Yk!ޠYdr0�v}��)��7]�N�}��2(�&��>�q���H/��V�!"}R�Zp�^ȇ�տ�A�uM��-@��z$�%��Wxׅ��ZJ?�=������oz�Za b\��ebbqD��tr�y�����}x�'�?G�?#TG�[�W06�Ԃk(D�w_ڕ��X�`���T�te�kh'��d�3��"�H���ۉ��:r���/���]��T^�sӫ@��)G�(�M��6�����f�0i�T���wI����e$�z�*�+F�!`a�p���b ����<��zr5�ӕ��h�c�N35��?��ؓO+Rx��I冻��KJ���Zc�ېG�F��8�g��%����X�o�ӗ+�G��,9ľ/n���O�-�H ?1y��V��5�ǃ��RAE�r"xU�8���(�� �C�twӏ<sڲ�?[B8�D�|���a�y��OT�8!"���FFM/[/֜7܇0{s��|n�u���ݦK/�����v�h�Jܑ�崤�j��n��h�?���a�}��P��]�&N^�U�f��!\�pd]�]+�Χ�i�^^H���d��Ӫ0P�V������^t�~��2XQ�x�J�.��kިi5�/�G�E@�ӱo�,ԩ.P��-T�y�ęa��F�!�~�*�|4N�Z.�g ���/9^J�>�:Z@�U�k�S��Ų��RF�3�KѦx'�h�Ր�0�cQ�u�/�@���r�tѦ���PN�G��P��l���?���\�Na5Ov�:�I)"��Հ�}��qA���C�͝�ݬ�_�L�\�L����,7�_��v�"�jxOE7N�8�a/SZ�a��v!<��e��a9��/h5�bZ#23B�2�{Q�XӾ��T�ߊ���q��%�[����a�ձ���=�0O���T�2�+P���X�Sa #R����y�ҵDi�KL�;�PQ�By���t�A�5�-�?T�faX㥁�F4���z��Sd�:�*Ky�1��Ț�&=�-�����gJt�,�:�`z�L�v�L;�p��Zr���LD3���8P*�oR{m�X�Dni�^:iE�3+����(	����~��{����� �b������PP��ݭ��B�q����7�����^��_h�T�Z$oxӀ���.�~mBP����
�,�����Z�g�oY@�CO|�s��l
�j���LB�+&CkCuwj9N"���D��������U<��;׈n�*8��P�C����,'�w�;1S0�U=�w�|b��- �}�Z$V����1I^_���*����"�q}�a�Q��b��n�_�~�I\���o���('�42���;�m�FZ�_�ADz1s+(��7�
�ah!��d��n���p�{�v��?Y�C�S�Nj��d��:@�v	Fp3A(7�\)��ؐ��L����s����g_wn��4�=�4���ZDt[6'�}�� �3=�k��SoWu!o���&��X�l>��w�#5=����Yv�a��5�ʪhpĲ)��9	h@!�za�x�B�x�&
j\�`
�!|ŗ�/�ku7B��9��\��Ⱐ����O���cY�de{\�}�f:cmao<5��M��Wz<�m������Ka����Tb���2?6�
1c�c�o%/(�.3ig����Bj�����dqR�~��k��.i7��ּ%��"�h2'X{	רP	��1˳�I}��t^��e7��6^�Y��v<���,�Z
_�c㌗=LR9��pz����3��pa�)���b��.��5W��@R�\á�������䪲ȴE���,wy�7�������O�4E�b��k-��R��<tʨO��%���GX��lm䀱��ۍS�iL�WA�/Z�W��R?/9��n��>{��gg���/~+�.��r�?�{��8ŭ/ɲV%Ӱ�g]�~t���&^䎞����d����?���0����ˠ���/�����3�)�\�${DHou��g�:P�A���1�C�'�+��,�G�`��P�0�	�yA(�õ>�D�m����'ȓ=dy�4/� rTE�Nh��D���/R��x��q9r#?-T�/1�,�Q���m5�4��J�>t�oY<'_	hŬ�M���7�ó��"�#0�d)y\�L�Vr�ppl�|<��dY�K��h�o�N|�3N�dx���y��j�Y͓e�3����ILB�R$�G���`���nU�k@�1�Wz�{�1��k��Ð��>�*!Q�/KE5�B�e1gI�G�:du�) i䝑FM���+��2���{W��a� uZ5r��iH�'���;L��w��~O���qC@R��E&��vKZ�@g"dr�?=�t�� Ԙ���P������B�`$�!�#��L0��4n��D�%�&����`,��;�����5���"A�;kjQE�r���I%���jj�L�&��F��f���%T��ک`�rC/�*m?q����;�F ǩ�Jcϰ�EXH��r�.uȱQ��u ���v������˿mp�]����ƽ6���#/��v#�"-�Pj�e�U^K�B�]Qj��&Gd|9��~�$O��_: ��� ݜ�X~�r��K{����XJެ�9�~��L��G ��BG�{��x��螎�H\��P�fЦuy�W�B%K���6��Uv$m��I�*2�Y�:���T8�g�K��G��)��0�����D�	K�4[Ev>� ��;�G�4�}�������o�k���X�k�XZ��r���=�p4��@���.�y�!�r�z]�D�L7bAR���
�-v���-�D�G��g���G���D
��g�v���9�G2����ᔔ�=oa3
�LV_��n����IJ�nZ�P�	J�(��W�Ut��
���M)}�8����F?-����>�sZsĽI��L��펟x���J�N�b�T�
H�#���%$�\��Ű�u�#_b+���2s���9
#����L�ڿ[D�E�|yp8�t��a�Ě	��?�����b0j$��k	��ܩF�+��;lRP9Z�]:r�X:r߮q�㤫'~�qB[�ꐮz햱��
z69�Pfy�ȏ-g�<� ��o�C�`�%nN��x�ϋ�C �Da�c�����/�ȑ���oF��!�C���ٸ�j���RT)q�b��5gu�?�=�D6����:���R/�װV�m�)�'XYs-��,��7ve&��7x�w]_;˲�:=|�0�܋�k@�'<��!��z�-(L��.+sy�!Ѯ%XN��ς����cǙ ��-]&����w��>;��j�ϕ���!(.�>W_�W3��f�f4�z
�T���RA Y�����8���^�����R�!����T�zs��?������Ck/Gɠ�rn=��D�{���-�|�sf�Ç[��<E��i�]��GmCO6����y���t��`7'��^�7�R���s�/����:��Q��&���Rg�D�<T�H0��Bz���y7��Nx;�[FK�>ѱ�u�R^�G�K�j�H��J���r���%�����LL*i?V�����"5$�R�F���]���&���#O��v� UG��hО?�?�]�g;C�e<L��캆7qZ�����ϡ�������@������̶�v��(�==�'M����T�=��c�k�ŝ���>�8颣����_k ����<�W�2��,ݳ��0e1��}P��������^�`�8�wD�9(��\�h�l<�YM���b������(r?���<���K�=�W�eW6c&b����``LrG�D3�u	ň�X�ӆ���"�O����}��7�C�����U/�Tj��V ���e��!@��ܣ��N�C����Ԍ	�S� �q(]�y�&�⫨��iH�MWJ��z�Q&P�/�ޟ	Ħ��T���(�l�\{DS:���\�c �L�:���B��=q��b�F����<�S�f��8���id�=��k����&׳>B�/�i��A0ĆS7v��o���Nt25^*�nذ�|��}�Z���t��mz\��9J`	o㬤�
C�N�ݝiKH�`�߾{��#�о!:����O5��?�q�������K�8��t��N2��W�uH�˪44�h�]�cl�1��f t,Rf!�u�ٌ{�焴�įu8TH��+a|�N��7�c`5k
y��W�ȳ�6�T&�}3�>���2J%c��Z�^ ��C���4���f�,�[�7[�xo�q�j����w�o`o��b8أ��y��S��UEb�j�k��T��^j
m�n/��
y��C��0LU��xWPϜGc��4��R_�����$ � {�ގ�FB��F<�wx���d�!χ�'�Q��.������R6kP�<��n,Q�\@�O��@Wj{AN}ɴ�'�s ������7R�,����O�o�X���B)H�+�}OsT8���'����uъ�36�C�G����lzoHx�PI.��G�j�uazw� ѱq��(��]���]�V��;Y9��p���۔�^q��҃"���y�zb�ہZKЧ�S��[�%4��RwM�J>D5?TǄ�/��i9%�\у��,B���( ���i�_�<,�Y��m�&�nT�yV�Wzs�I�J�, -�  �>:��ʿ]���8�F�5���r�V�N���>�ahhZP(�PU�*t����F��$��1�z�xm:B|'4���r/�9HK�,!}�Oɥ
`�ꍜ'd%��3/��p\U���+2�2����H�Ԩ���xv�͉�2;�D��uc]�WZ/T�f?�Ҽg.p+Or�#�����gSg���+pҝ��(F����<��[:W�VQSu����N���I��	V�lSuf�>:�p1_�Y�U�� �l[J������	�3W�B�+��x�(�I�?�O��L����n?��J�؏e��X��6{�L޽A""E|�I���ٰE�D��Wb���W�A8]�o�]~�VuF#zE�6���,o�B�1l1)��jK��Ӑj���1�(��n��1�}E˗c ��#^x�@����3H�5/�E���-��KW��*C�}�Q��~Q�Ʒ&vE��~=�7��x�#��d��j�"��I&�p\q�u�?����6�4�Xh�ɺ��Ϡ�B��c��,�P����A�~O����Hnf��i4�~5�:)��Y`0+�t(��Y ��ձzp�C
u�ca�4NK���Y��C��6��Ɵ(iC�BǁOgU&h<�L�4��;a3�^`u���R#*��#�>|��O�%ަG}�m}�1�l��!���K4�_��U��՟$BKLT<L���C�p�i���ұU���So/��^BG�G�����A��F�����4��c�cz{n�:R�)���o}fx���%Y���e��Jkj\4�c��&���1H�
uq d)<� ��'m֥���Ǹ?� k��y��&s���]-�$�&qu��F:�?A,:���l���ҧǒUా$S��C�,7�g��`VE�Iҭ�:�k	��Z�����>��k�Fb��)�ُa�d#������4`����%V��%~����STFE�"��ːb=�]5W�%�FO����t3C�����(^fFV��HAW�4���y'�/W��ۻʒ�$: 7�K���baڂ��GQX�"�;f]ٔ�1���Xk��ܡ 6^�pN+n�W�cX�̓j��,j��k:����v����A�4#&����u�{!8a
+�Y�Ah�y��)!����-.����Jq�t����N\I�Uf�����_f�S� =��J1�#��O"���ѭ�V9Db�䖡��ڠ.CIS�pC�<�e[?�V�4R�ܨH�s���X�*U�H��LY�	U����`�v�7+/�b~�W���i����g�5΃��A��f�ͮ^�X���բue�׭�Չ/�.����G�K�w������[�[��F�s8�{t�15��yGNL�Ƀ�`>�Rc�j�����&��Qo����A&�IX�nvM=� "��t,�������^��L��G�q
��rfV ���J ��`"p����Á:�"�0$� =[/�B� ��{8�x���	xQw�\|��� �=��
���m˃�;,�D!���M
إg�s �J)2ͬ�\�����HJ/q����4����^��I(E�	 De*���,u�}�3o�}ər�Rr���dRY�0?g�YQ�Vre��.�v��+;�Z�R���� ����+��6Vj�_j��Nq��ȓy�״��n>�K_J�9�F�k"S8�M�%`l���e�<��Z��|n��R>��(~�W)�D�>����WX�%r������M���YI��
���k$^4׊ۼtH�q��@�Ϯ���"48m�%!!�R��Q��T{4��������}O�e���;��a�=��T1'�ܙ�q�	Kr̻��'��������)�Y	�[{̃@?LN���8s��/�F+��߇b�5���g��Da��!@$�h1��|�׫j�(t8�,�i���18��ހ���c�:�lq��gRj�~Z3�L'�v���}K�rA���hC1 �)fw�
�h5�%#�B�
�/�j{��#��!��!��4
F���F9Z!�3�e2��p{�0/��>}�\�Y���T +�C�AF��vNQɝX���#PSPVk�@��ߡ�U��\�Mu�Y[�����h���he��&������A��ƛ��lyr,�����$\��8�������õz�Wv*��Ra4���}�Ѥ#�f,E���pG��(ħ��y*�����M(�a��k�otq�s�k�W��Nĳ^s
��ٰ���v�6*Ǒ�޺��q�J�s�J��a#�V�>�C�7�K��o �z���eJ,�e
�ύ{`�8��EK�&�nmr^<mAW���UA:�b�G��`��������n�na�������{܇!�	���Ԧp�|3r�%gf�1sb���TMë�R���VZ#,?콥9G#8����1͋ mB���˥�J����	;���Н�����$�a�6j.B|�t^�+P�l�O�u�����m�aK�~�A.��bh��7l&$�zv3{�9E�#����7���#��f���84%y�(z����>&�������,��Q�����7�:��_�DT����X��{�.B���8l��,� ˂ì]��)2��g?]_ �C&4�+%�h�;@vs��<F�uo۩Ǩ#I�c�]�;PDU�j�iK#Ms���tf��3�\_H�����38�$�sεN!�ݓ߄+�y�.�˽�Ll{tJ�Ц��6��u�8�g�iU�QZ��F�������K+���#]�}Xk8�[ƴ��No�o9��?
ܩ�/2*�>��MK�C�Ժ��Ox��꓅�e�QѰ�ܣV��~�%xϽ���N�g�L�ⰞhL#��`�G�Y]�x�*oDH���3`��t<��,���'3��
9����%�}jw=�Op�.H���G��ܚ�WF�Y��O/�mv��H��y�_�E�ĉ������U�[G�+5�%�̔����[��NO�^e��`�#�j�_j�I���O�C�g�e�c">��tK�1�]�l��IA81Ĝ���j��)�-�Q0y�>��)����X�6*z��:����`�y�舓:����R�$�~�����{�B5r=���ch��V5rv�^zQ�4��[m�f7H��v�7�DS3w�2f��M(*`��+��c�
��4[a<ϖ�r����(�A�}�@�X�.���[�.��L���^K�P��L;M���y]G���0�.	ۡ�p��J3�P��D�l2J::�ǟ
���2��5.K%�0ަ�i��#Cc�%�`�����?�	T0^H_��-��]E7�S��@�V��������t�R~O�scDd9zI�J��3�^��	$�[ް�_E^,�S�[���wf���8���w� �k-9���c�z��+\���e�P��+I������}_�m�r�:�1y4�W�>�G%�8�d�M���\���u��;&ͬ+%��q��f��<&����k��j���E i��'5P6��3�"vB��ZB�����?�)�N7p�����g5+���nt�s[
�-����n��&yUdA�OR���`/&�2�	3�L���{�F��F���O΃=Nd_�����H5�d�dw����E��9"����y`�y"�ƺJsp�&����u����$W;7�[�3���=�dw�d�X�����8���-c*İ7Y�n��w.��g�}��A�8R\H�E����ˢq;��ؿ|��nO�%$��z�@G5H�y]1���q������q�����z�<<v�}�۔<�����:�����^��(�Q,��g����H�k�
�PT����[��z�Q�_��}��E���D�Ak6WTX��pm�i*#�e�������Nw����-�'��<Q93" ��q=�(~�n2ʯKZ���o�X#�g�n�A�v�M�t� �TX�����#ˇQS�͎B���n'/_�ٴeִ�"i���b#Q�����-9.��"������0J;�aE�&�%�)m?��7��tdC²J�ùI���g���P�瓝'O>�����:`�s��U�j89�A:��ke@��Q!�����q���@�ml
Tm�xc���R�ґ�B�m�Tva�&��'�,�ˤ�e.�h�@���x���O���+���Ό�3��<�t4X��Q�38"�������K�O5�U�>H�U������-���'��Ա�sn��[��� $n���#�H�%�﷥����o0.;ߛ��kQ��ّ��>P4�4�)�Q�<\�Dyh@����ΦN�@��J`w�ԃ%�ថ�&9[k�wt��G���I��/���ڵ�A�Tx�ڥN�7%-��b�ƶCP���������̯���ڐښWt�[}�el�R����j`�v�k"#�Ә�Z��jO$j���	�n.�[ϑ�s��vgZũ�|����ӯ��Rݩ;�ſ���]0��wU�˲d�����J`��-5 îJ�r%<ɕs����A`��s+�%��$�L��yZӪ�������Q�����:#�^+R�bH��_H�@�%�3����X)������o�`:�cl��,� ��y
�oK�c���Xա��5�[�sf� /f�,����8d���r/���D�7�B��㼁�if�́�~䤆*����87���09Ϲ������)�w�߀�}�z��&B걂��-'5�~�7ڈ	���|��e(���������
j��,�O~�~{�`��$[�<4�>���}�y�kq���ḥdh����M������\�Z��o��G��� s٩�3�"w3�&]�sW�j�P������6��h����1�m(�.@гf i��=����~0�G���4\�d�|F~���
�T˙5��}&v	��xb���J�X��>�/E��P�3�- �*��Կ����?�K֮�ej8��Ւ
�+���t�y~�R��Y}�z[i��CY߆G��)�{4$�U2�v,͢(7��!�6���WR�$D�v	�[Rz�T��Aׅ����:.swZ�ss)fT ��+ʿ�\O�S]zַk���0 V�,q�[!J*���m?�:�:>7/��Rb�0�;����U}�F��gC�1;���B`(��4��H��mUt��#�c���+Hs/D��9\�,��t|ӳ#T��^9Y�_Y*.��YD8�UM�ޏ0N��D��r�"����4�`X7v�g�B��e\���M_+m@�<Qg!^���!����+Ơ�gA$�/�Rx�q�K����������Y��8�6�մB�U�t@@�~��J�F=;��o04}v��CG�^�� X�4��0��隢�k�9($pd*x��F�U4������8i*w��G�S���V�o�����2���B��6�k�M��)�����\�V����k�W�4��m!��K1[�}�5�t��A*�t'��[Z��9Fy�ڑ�u�a?����J��a�J�0iBF2׾�J�|]"���R�7v���@w�B�yc=�c�oaIʂz��}c$*���uh�<jfk�9T���\�YvZ�J���G콡&�p/O�t�/ڲ�x���,̃���?c9tB�f��b�}t{[SE���򛃂{�"��m�i;�ļ��(��R!V_�V۱D
Ԓ�ԕ�#��N������VahS��Y;3���u��� Ҩ�I'O���@|=�H��}���+b�����L�d�]#wd���_5�l�_�%�5���D3BK?v�N��~u�q
�!��gU�4r�{��gj��ܔ��X�ڑY[���Ѽ6����ۈ�dT[Fx�>���ϸ}O�o`գqb�YB���[�Ӄ̣������7m�TQي���Os��K7l��p�F<�jb��g?��t������(�6y;�Q�v��G�K�HT�{�����_�[�q�+i��΅���ؕ�+X�=��Gy+PK:�����S���IK����50�ť�:�!sP[�* �0���Lp�Gb�� ��Zְ�����7��1jy�&a#�Gk_�:�p�cM���IX��;*2��_#��f�����+/�)qIW8�$�_6��������H��x���A-�hfU�L"8�Ƙ,�|�J�A�3U!F�!�GБ�!�S��`�i��f�3����h�*݋���˟	�E�a���,ժi��ǯ��� ��r��g�����c��v��ꐜ�2D����_]��y��mcX��Fx�-���"��/r��!e��0��X̻,��������w����q�3�Z9WΚ�\.�V8�6�P8 �[����/�*c�=+	(�n'8�|U����bw����]��u"����"y�Gv3�=_�䎰a���{��&�lx�q����q���uJw���v����������Mۀ����;���������ǒ't�uǀw�,x��p�d����,�ta`��А�湯a�5	�>����_�L���.ߚz�o����}�[x|#!��J�'m�,4`�ˆ&�����
R�n�q=A����Q��C)��6I�v�|_�Tn�;�FW�J1[��VK�_I�-�Ä��ub��}�Fl�Y���)�]ș���/������ n�t��z��Ӑ�#������u�����,H�/�)�Nբ[���`nR0�'S$f��m�Ju�8�"�L�|"�ޞ�S�7h�#�^Z=s(ㄋ��<i%?p$Q�(�Ol|�I$c�����	_���
��Ӧ�:�(�va�{
[�h��@X�m6v�Lcw�~J���4����N^������l�Su�����i'�±i�Ѓ64F�D���׭a�@���/�<�s1����Ɗ,�|�� 3�|�]�yTǈG�]�O�aN��՜��=��d�o�$�l��
���sTh{/��Sʷ�t�)��T�A}�S5�D��BE\4F�*������ލ we#ʊ;uZ��gHZ�Nr���F��9I��b�bYUB�^��Q��J�t2Gh���PX��m��h���^+��н��2��I�t�Ynob�
آ.��0yh�m��1��aFfc�ʈ���ˠ����o�~6�e*�b�9�-��E�=L�b��	�ʈ�ю8���v�5��	�0ţ�fЯ�(��eK���� ��>Bʁ���o����&�G���4�b��+�[TuF����E�W����jX �)�N�����gq�Ţ\��	;d�����=�`�E�B�q�<9��?׻�����;��&�UF��ԭ���ǲ��g�݃,��~�~C��I��t��b/�v��Gؿ��t����Ĥ��}���u����˻bs.�{g�躅�h]S�.��G��BM̮Z�]�^}S״��b<kẻ9B�Z��$؆��B���daTAO��c�:r(��|>s�D��L^\���g�?���-��g�-G�����ImW��LT1HE%��txr�[~W�3�n*Γ�'��K��O'��0����6<��[��iN�WTJ�hI�K�ЊQ��VR�{
�=���[��Y簑�[�5��3��&�F�z7��;4v���͋!����8�Tf��u�����݋ݸ�5�F%��=hm�<C�Bp�9Vq�nˤ�w�^M�m��G���( �(�~��ۛF�����-�e�����"v��tr�2/d�OCU?�Z��tc���E0���8����&��'��L�s�Qx� ��JuG�B ]�~D���!�r	1��"cT)�gO���T�w�T�������k(���B�z�n��.����G�y���rݠ�إ�&�'�玠�TV�09�k�ڥ�� ���k�K���(�z�T�\ImWq@ٸb.1R���ȃ��W�P^B�H��ۏ޷��I24�����|ǆgi%�U�����j(����l�,/�j�;����IR�Ky=4\Yr�Xt
,�'���A���
	�]�6 �x�]��kl8�@�S4 ��'[����N9��\	��✱,�%O4��	 W��=�T��"z��u>Ta���E�1Ѻ�pJ4��}?��1F�*'�h��L�� +��
�),A&�}C�Jd�K�0��n����2�(��-S���n"%[�����!d):[���A����q]ޖ/������=\�`����@����i�k�~ɲy��r�"��#����޹��8��Ԙ6��X� ��Z�A�^N-�
,�^��%f��t�$N�j���><������6�hXu����_p��"V�`Љn���)u��
� dK߷��%�##�����J̒�KN6�����ԋ�')��N\ufr�L�%�'� q��
ºc�W����gNAy��)
����q��]�j+�#T�����C��L{�+鱜���Jz� ��[Z�k \��P�/a�a*�B����~�V;��&�+L�\|[�?÷gb�V!g��$�y"�;.p�����)x��Lb0�1�N$<��:c�8��|Jn�m���U��c��{��n\���L]�#��E�GB������Β�����T�!�W�L�i�
T>ZUi[?�P����c��Q!�3`ܤg��V�#9�A��4���>�貁c�70�C�{V�R�9������m7���@�5�i�_����ż��T0^z��3�-L������B��Mٳ�S�)�%]�ZkV�a#�U�8��"й)�4ߤ�2����x)�����j�{�������Cv��#uX�b��M�-�C��n����:������RA�k&�b����!~�G�JD����z�nGF���8��`鴆ܦ�۵@C�9b8��Ls�*z�Q,�%�{��g(X��gc���
� �@���У��Ѽ�-r��	���f��*���������2��<�m|����57&H�oy����1�S8���#�ޅu)�[l	�������V��J�����[ߌx�$�]�ത�e���&x!b�ڗ�y���a3��Ss�Yq�w�����DY���2��C)���>�W��ȧ������^Eif�3�G��X�.��-�^
�<B'�
]�j��f?�ٟ9�$�5�He2�룕9�M�(o�v���L�U��h֩YW �27���0eA�}")�;gF,��i�f�|0�C�m�p�e�E�G}b NE��@��/0=^Y=c�:iWp�����K�,��ȃ��{������\r����`���	��k��cs�ω�e@�HC����M=��Y̚�h�YU�Cv�ZK�=�a�ћK˜b:3}�'Gϴ�[��Ď�T`�0>���B6)�5;�^��P�z?���5ɻ0uGJ�8Eٛ`�z��i��,���P�e87x?w%Q����y�����9���\�.L���9����h�ߣj5j��?qL��@KJ�����p� S�����[����6���}j�Ѵ��Uo#��!�?��Ch�XJ�rSz<�o�H�Q�$���(}MDP�D>u^N���*|���k\���O��i��l��}�_Ieu�~�3@u��j�]`��F��`a�:�2���9y
����~�R�[�ͷ��D��H�k
2]�q(�X3֯�Q�� ���٢��@j�.�l����� 7i�G�-�X/�K!\�C��3BmS�v��m ���d�����?>��gjU���2K^�#*Ҁ^�qG�D���\gk�d�����p���T��ZP����'�d��#�=���wSw����S�1�
�hNi��ÍA��Qr�Y��hi�+�y���qn�/X���Sw�>Ċ��
m}�^CJ�f��/�[�e���q�W$B��`�����V��>zQ������>�I��+O!��`g��*�����=
g�c�.�*Ҝ�-f�MM���Ahe��*��z�-���c�ݚ�x���گ�dI��M�	u�
�1�����fȞ�)�t��l��x)���H��G�� �*&2�� ��i���a��O�xݵ��D�a�qʝ�$�|j`��@M($�c,|ue��{�#�FEA�t��}Br��h��� �ZF��|H#�ブF؝�c�K-r�N<��i>�J�+�OB�f'o4�����}�)���S*�.�'����V��٪��у�+�"��e]=`�w���"M��`*� �d"t9Px��;�7��ײ���Lm�p#�v��	�{b3cIaL�T㔒WL��0Đ2��6_���͢�����w���Yd�I��\WN/�$}q�[t_~5OĽ��B���!�ٕ����Gi2�On��0�]0���JuD	(�ә^2�֣]����lD[��H��2w��U�rN>���:
!�{0��ג�����A�}Q4��N��*�x҂�7��Z؟)����1-H��߾�"b��?Q�\բf�gz��x4��dk9L+�ֻ�Rm���6=���,������zb[�q��ۣ�Q�t�Ҁ	A�g]���{�I�k�:�i��Q�U�;!���!��@R\��+ �ښm���J.%Z��%I[䈩f�R��0 d.�%ybĆP�z�Ni��A8��'E�-�ۿ+U�}��]�m]���Y��f*�YiU��vl>� �	=���Kj���La\4�dYQmљf��Sut34Q�U�(�X�T��~��HY棣�Q�4�i�C8��a�n��L��	-
��lVf'�\��`r���2ᢪ���\��a�H�/�~�����n����حx���6�ҳ�,X3�`V�ڟ���3*�""*J?���Hd���߀K̙��`G��z�g������2HƗ�_��u�u6��
)$��[۔��U�VG\�Jq�B�L
A!��n��j��7i��urqA�3Ȃ�6�0�y�~Ӫ$C�}�G
�6�P ���n&Ҳ�b����w�*�� ��A�7w�0��5$ ��M�}�����yx��������=
҃� ��������d>[��zM�~�-;!���'�/�P�p�Y���!��H��n�|�|c>�'��p"�9��6۷@��1���X�m���	�������J?�����{��ퟕ9���/lx)�,sq�ҥ�x��|�~%�΀q: ���C��	��S�V�a�ENU�c��Z�����j�n�w�^�!D]m-K澯f�B^a{C��� �Hy��^�F������?Dͺc0 0����~�?Ѳh�%R*�dVU�pF"�7���В�Zp��V�]�]翝,��V�©mʄNP}�#��EoX���|=Gk�n�'_0_�kTӐ�;a#��Yw�&�A23i'�r9q��S�'�2
��A!��9Y<��ί�-�E��||t��k>]K�ܯ�F�� e'�����^��F{:�k��h�A_�h��n���e���?Z�2�2Sc�;��e�7�T��'�H'w��% B�Y��N�X���Jq5��`��D�!�=����v���R�y�ܨ����1~ƛ��;6���&�[�Lo?�i
����a�T�1�����Hjr�>|�p$6^E�l��q�̴��|�{U�>��ŹNg��鄩jOd ~[�^�Ei��t)f&n�1פ��ң�h���S�\W>��"\�ʘ��<%���nTT6�����k[>�!J|(���������:t�ڣo�y��=��ި��F�=>���A>�O����*	B�H���
��Ȅ�^��i3`�fz~HV:�S��N���T?8O������#b���"��z���|�h<7x���#���3jΗ�v*�	��<5���7T�b:��m�\
:�es,%����& 9�D{%H���@��P��[qꣴ�$��[�Z�[H<�Y�_P�����Q���ZW!�ۖ��B)l�3_��zM8��7�qʵk�2C���o�x�f��!��"���cY,��bɚ4�@QXwC
��/ ���>M}�CpqO�U~|�����:�ݐ�ג�dc©�|�~ŗ�����'�c�ۍ〣��
��͗�G�.	�7焐�C"�L��A�OK^	ErSe��G��$\L�C��@��QG��VuĠI�f	JW"��[�y����7i�o�򪾻�1'��*��3�6Q�6fZ��a�#Jf"���h��eOX+���p
����i�-g�<❫�=�YDo|Y\���� ف�C�d��7xU4p���}8!z��;Wf.�>ÇpmR��s!����+u��Xmɫ�/`�M����ȶjT-��m$*y��k���2�f�QQ�LK���w���(���T��<=�v���wW��9���sH�(�#��XH��1�ٷ!{�0�i�>K9���L=��wF~�T��������sA%8�m��<[-TL�z54���\�a�w�`��Kq����"n����ʘȕo��1��{'1�����I��l��`��q�1x�
Y�틏�s'�f�T�e/�4�%h@7eB�aJX>�GDO��A�}���P�;P���K�M@���LX��>k�� ����2E��l�0d��!��}J/M'�4z�\~�z�z5ol
S�M��r���!3X�B�U�ݩ�����&��,�9���m.<B��.�;��	���p&�I�jA��'�J�i���؍`!����(]�L�t�|��S#l��T��������g�QmL]٢�Ĕ��ɋ[���%]��Ĺ��z����HԠ���V-ܬ
�{�����YwN�?{⿣��KD4x� M���^�`�<���;'jy�+~}rژ�ia���x\Y�^�#��C_�=�m�������S"R��H�~�����@���=�ē�夎�����q���)��(z�K��6Ԍ��D�b��Ą:�.Щ�Y6!�r�U����v��j��{�ȝ�O�N'�+��qkZ���u&]u2������󤓜`"*}�j*a8��N~E�4�G?�ޝ�v���0^�p���KЫ������"���g8;���9����=���I~G�_�KGI���A2�zjoud4ɐ�w]���B�v�g���wx֖��F��T��X�"�7ί��o���L?� V�}��j"s�a��6Q�UtHX���z�)(�������/��%j;�UÐM��ǔ�v��Y��8,t�T�΃���_K�\s��!6Gh!��{�@Ӣ	kԽhX	!��1��N�F"�w�M��v�<��猚-9d�m=y�syWɗw�����p���P�e��<���v|�t{gf)�S��-���'h}u-�G��ՙu8��^Rv~a�oe�q�4@�#I!�՗$,��A�!�E �7#�C��+����m�zPQ�~v��<<k�:E^���v�m���]_+���v�#r���x�'�S��O��G.�p@n�F��m�&	}!��q��CM�#�󑀆��{y��#'4�8B��pǶ�]?�gA���3T�暖���G#��%�U�)������S��� x_?���wL�2�di�:�v~|��<g��dL60pBR�}R�`��.)��>G�i`յ�N*�Jj2�ɋyv���>.IGW�(#�]��5�*��.r�M�,4����[Ʈ�n_�S(��J$;A�e� !����p�>�
��=S�|���X
��9���-"�+4�k�"m}IAт��l�'�貦8X�hQNq�<�OZܨ,�д���������[�*��C��M���
0���W���l�dL��?]O����Bd$�l�a��#�4�Z�k���"���۹AY�^�Q���-�_S�u�}P�$�����,f�}�s5�4t^	ק���R��m$��rR��<�d�A����=�x��Vj�&2i��˽cɌn�ª�F3���vB\���85�,��2�^(l�-�� �n��ك#�Ph��J��O�[b�DLFa̅-�M��)��Ǚc�-=�(�Ly��k��.���M����q����(���c����>�|�ࢦ1�W�;Z>g���ӂ3�w%`H�w�?xȼy���Qw4h��T�ΑBƵ.�����g+�+g��Z����PU0YR��' ab����q������0Gۙs_FFi
�IkП����J�-�z�yfn�Ն��c��P�|f��4m�f��X����
{��~����7B���@����hpn:*쭿�&��7_j�ŀ}>���r\�)�\��%����B�D]�?��r�x�$i��QO�h�;�6�r[]6p@���2� c{217)�cs�à�Sn�W�sDu,��g<��o�܂����o6�~ʭ�r�X�� <=����s�׫%+�VW��"<*���e+R��xN��	F�<ҏ%�lӧu5|B����B���i\�=WaI�0�2y��!�I-��53��T�u�
�;Zr|(uՏ��$f���YL66׷���仯�E�d�r�7@�g	bx@��(?{�^L<*�wO�b�{��6�&cB9}���[f��<i?�H��w���\��N����0�S!M�-��ߦ^���_o߶V$��wvy^h�!�m���d���F�N!��G��כ�4�����B7tΎP+��LQi���ڭ � �M���nb��ɽ�߈G������4=����n6�]u�i �#n��5�G"��JF����>�t����0���^�leԌ�1�;8��������1���T.���O2�����`]����� 뎱Ў#w��ރh+�<���L ���rW��tM���X$����;_B�z� ϋP~�t��
'�F�OK��>��󱝯bY~� *4��q�LQ18?�^W�%P�@+*kN���L<�< c����C���.�-�2=�&�Q�mɶ�cq\��!�=+�cr�����=G�>�f�%Hms��<�Rwu�_�]�S��"��֎}��:� $@y�C�n���?v���(�,�8�YE��������0�Wd�EcK̉���&����0/�G*n�*OY�<��?��B�Ͻ�BI���#XN�q�6��q@M����[jU��vpۗy�Ki}=�f+�R����,I���M�^Ru�hgQ�B>�֤wU'�iB��{�d�E���Yɓ�S�rn/@�^~�d�n��3� �Pt{T�3�����b��|���	���ޟ�o��G�����u��ED` }}W���zt��6d��@xkty��&2v@aI�	ܪ�)��d�L9�D����Q���p�4�$1���d�Pb�PLd}w����t/�7L#���9V,(�'����N�r3��@���aԒx��8oo��l��SVa�z��Y©g���2�����̨��P?�B1��7ż�ALw��)3����l3�%(�9�=+8,�M�l�D0�h��3t���U���b��U,����R�h�̅��(�F6w	�A�@����SŶ^����^���$��C����O��0u�(�Z�'�FY�)�|�V:J��E������f��m>E#� n��I�o�䅉��,��k)�]����u��{-�O^v3��>	��$a[J5&�)}F��=�M/�!�'_���E��Z�SE��̋f[�d��EDL� �V*�1�Td����{vқ���ڞ�5�Ү3�4ٽ-)��߱�(�j\�L8��5�1@�hV�}�m��+FK� ���������*�ꕲ��#E���WBI��u����Euh�%�T�j�7SުF�mɟv��Cmܨ�hm�Y�2s�俬??��Z "4
A�ś�Pr��yq,�{�Ҧf��Ã�]J�k�cÜ[�6����N+�N��F����XOy�	�G/�N�������"Ĕc�}��nc��7XnT�/\�'`]2��`,��~��ق���e�Z��YK)6.S���F��*�U>��Z�84��Y��/!c�����9w���E�8�*Ѵp��"�Y������Q�T�2~Y���'z��,@�[j&�H�'��SRM��K�ND~�&=hps���M���a�<�D��n�g$��R��Fc��S�����O̊���@�?Jzä�h_�	c���sܣM+���Zi��t0�5����:�'�/{v����N�B�$�%�|$��NQ��[�W���.�G�z{��٣C<P@��䐺'1�+{��V��Z�3k(�b����%Jt��	��G��%�v/T9L��&�"�O��,7*���p���<��Nc�W�0�>D�j��@���#�ĒJC3�޼�t��y`)��Wy3�O�VX�E�E�.a�\4z�]��V��:�O�Vu4�]<߰�BRbE`�݋Z��SUϾ���(F×u��쎋
u<��g��<at���)=b���j��}�ȟ�_��&�(��>�Y�1��Zy����hX�1�m�I��B��v�X���Cc�3�Z�=������#���y����W9=y��T����)�4j:��n�j&E�HZ��>�P{���g�,t	�Y����ĸ!P�ZyXC��ׇ��A	��N)�!�RA��i{�$�g�V�_Nh�v�=k��@({�I�87���.��`�,T��%�
���}\C�w�k�a�M��T<�m���a�8>/g 6Q	��2�\�L �j���c%�SD���#d��[�r���5�!d����BkG1PS��'�/�V�9�急��ZP��^�FXY"k�3C�uI�����4���D4����b�w�,�Tq|e>�.��-gG��uA4'~A_N\.�����dh����O�:�f-k�A����B�c�����e�9hl"���چ�F��U���̅�3Md���g`d�#b��=���;u3,��;�jf�(���%!����%⊜�.r�o
�5Y9�c��� �����*�̭��,+^��&���ť��{2B$qvz@cM�OU�q.�ĭ�F�\ap����V�02pw*u���q^���9N��+/��~Sܿ��&�l:&��&7EF�$4cao�h���5M�X�#T5�@\Ȗ~�܍�6��
���֛�'jn�O`@�ak�~#ϪmUD-A~b_[�He�;�E�K��"����Z���t���`���X`��aj�i�Y��Zs;�u�F��5�m-�F�c��̏�����q^�S7���03�ty�9o�:�z'QCG�N��ʹJu,�Η@�7C%<���X�d�d�]<#0hb�.#��*�@aW�Xe�1�/Ҟ���t4D�Z۷nS 5Xc��<~Uŭ�23ot%���Z��@Ҏau�M8O}���0�oߚ$�{������{u	ف~�T{xZ�S��mY�1���{�@�@��� �|�R��E�����H��512�e�j��{�Pg�R�k�*��70q#Z�s.J-�%-�z��~�$���@��e^��S�����a��%W�����B�e"�J����bR3�y�tѠ��+�2[f���Pu9KL���H>�&���N�y���Q\1}i3�4%����1�V6/��pt|�'����e�?Zȣ�44@�S�W�kU��x���`�XyB���?{�y<$#D&x*�4kN�:TR��!)V}W��t܌
Y>�c���02}����d٫: ���_��cBA�4cL�!u�J�g�+~��5�O�%�s�<�m9��Ʃ���D��?uaK����r��4kfp)����¿�8OS]��;�5�۟���:Vձ�L���A��J �'�>�c�S	W�����iݒ�������X2�_��U���#�5{��s��,����k!�8J+V��l��͸(M�ڇ����c�;��]��r���C׮v�;sȄ��hM �:dH9�����rPW"�2n���|�K20u������poa!�e�0[�z�#��;��w^�t�0������abͻFߊ1yW���nA:Z�?ֲ����i�� `\�� q��A��kj�6'}�W,���.��d��,��mW��R�M�<�u��;{6g�yC\��{+�|O�H�^N�/Q¾�� 9��\�s!m(yH�x=�Pw��Nn�����.�����V_���9��[��$I��iCa�6�UIB��ʪ$��{����թ[� Ҵ
#�b�����N�"���nc�8�T�\��yf�Dk0�¶�T8)p1p��o��0�^��?��P�EpK�f;1�s��#�2���K	6<���9x~�L��"Bm���+�MBn)����x������[y�=�~����g�PJR�Af�9#�=�	���4G$;R_���Og�d��<�'����&���$�!x?��6�!�~��oӝ��m)ǟ����>E�)�<Y���f�9fP 8�}�ƙ�7͍��Ͻ��K*�_���k�Wq}�<�N�ֲa֢�����ײ��l��䔖�o�c��c^RK\	 U]7���8�����1�Y,�*-Oa, �_Z�e��� �bZ7r� � �G>��q;����x�B�g���E�Z<��|<ט�.w^R�5�x뮁��BL��2�����Y��̗@*3\�$���F8� q��}LO(�)UA�>��F	�4��'`�@�dK/Zæ�aR�z�t�9Ot���b�lM�*W���R���c5|@{@��+IVQAkJ�������bm�Mv����I����<���ߓӛ��|�r|�a�vO���p��R��0���#ƫ����7��F�I�����0��Y���n�gyO���o35�f�6���������-!�����Ė�;C�<�n!�5!b>�/�����X�%i��0*�;�W�������H���r2w�fX�#7����\��.� ��jՑ���P�ɂ���4M�1e���0��S��\��U+�m�%&w�iyׄ���3,F�̇����\�G9�q�$T�R�Qڜ$3�X�id^ 5������*ݷy���@�2�p4�b���@����Ս�*'�O�Q�&T�qD;	�"A�u�"�g�'���8%���R�2�8�3VZ!��&z�IQQK��2�����#�<Ni�Mn���3xC(de� (U]�9��&T��� ��|�4ΓwS��U�vƠ��Y~F&A+��o	�#uҁ]�5����1�)y' �8)���5/�$x`�r3,�s�3������>!����5F*�������ܸm���B�ge�a/�S���K����@���E'''�uA���3_�L��Qd�aQ?lKD��e�����6e'z�I� ���A�	��!oi~?�O�j��y���iXP�P
hs�[���5�|3��H�H=i��̉�ٷ4j����AA�_Z��1'I#�|���=X��勬�݃*M��{��t�TQv��Jɾ�M=�k�>�v�>/���s2呫{�Q�s%��<Xʄ8�s`7%�9Xa:�F	x�H����DK͔ ���	�x8�1��Q[�б��b��wȫ��y��([�f�6��`yVN����|,��WF{tj��:��<����Y%f��dR�J7	XV�"&x�@fd����D��oҖ^S���@Ra���H�yl����يK�(џ·��L�ɤ��["!�E Eu+� ��������H���;�W|�0RT�k�&7/*��Q��[K���F����G8� 2ow��	�� �Z�]lЃ_�X�T��^�v�q��_��V�lxt�g����25�y̆�VF�jW��~�3�/�u���|[#3���*���� �h;��K6�P./`GV�c���l̞�W�����d���.hT|v*��g�Ӧ��?��D����'�ھ��1D]��v-��かe<5��)\��ˇb*�|1�<w�U�^\f��f�]������Ұ"��.���B=[�Bl���<���lDt��~ԯ /��jc��h�Zǥ�YV�_�y��5J$>��p��SQD�s~4	%t}�?�P��p�HTc����Uf��t3�JvH�a��Ƕ�GV��߲�����`U/��jf��[��U�����@2E�=,]{��,�3�\��M�G;��̶�^J@$����eO��r�M��������Υ�ْV�k���z��3)�[~K��n�HmM��z�4
Z�ګAq@���"�FB���� ʕ�<��39������R!�o�0:̭$�?�T�^�n�1I���@"}9D�9�r3E�����g	�Ɯ��9#~�Pd�ۼ>���R�j�K$��ߒ+߈���6#�� �"q<�(�uu?�	7�(�=�]҃����W��ӗǊK�MK����eT˪J�(K�W�!�R�<ӗ\�?�pFudUsAH	�]����;Ɇ�h� k�R?	g�H4����p�݌�� ��=���0gt��).�<ԡ8���0��w��8\���%O0/)�E�~f+��-d�Û-���3��;�[��I3��nxJ�I2�`�-��������d�s31�;�2���CTy�Wz��w��+�j
���F��x^�ӷz�աlN��+��p�����V�
m���Q���U�-�E*�$�T����w���������)�s�o��G�}�+���H�sV]���A�y!u�=T �cB:�����~=�Pgx���_���C� .�$a����X�3���{�t� �є����%�Aa&�MP���\���S���s��E\.��Ü��4�m�V@��}�	��>9��y��?�G�D�~N^�R�&)�	��s����/f}���/,+��ӧG����H��ˠnާ@��	��ٶ��0�qEw8��v�G;?k/ǧ�Q�j#�����)hvE�7��{�})�lc��Q�S${:�-�Oz�<��q;�����f�)C/�0T.�
6��o�L�Ȇ�'`� ^Vs��Q(��"s�o4O�<'����D�h7�|xraL����&j"Ή�5�1�����b�y4�io�ͧٸ0/
�Z|e3�őL��9Vu�-�WH��$��7
�:F��(���k̂������(��|�V�?�Rbu��Y���G>z�Zo���z(���:5t�1�3*��e��7NĜu`x�̹�1둗����1H}u*�,a&S��t�VtN��QGc���G�v��|U�)�d+c󺬶���!��=-�!:eW���@t�T.roS)���]�ݙ���`Ew���>�P��u��ɒRń�p\&�����f�zt��������� =�iY+���R+�0='��FG�� v�含�/��P��<��[3|�U��/�,dVq��<?2=��Ĉ��3��ba�"/�q�QPH�]����g�6G:��a�	��Y	bp[��Y���f0c�k�S�M��15��bt#d����=.����.�2���,���}�kw�x���
��n.��]���"*�T27�qп��P����Y��t�-;k�N����&~/���$h�#�x��u	4U.d����S���!���3,�?�)����GJC�!C�/�ϡ���.8�?�Z�!q㳤/c��q��G�
���N�0!����\�B���o�^�M���(�q	�f�*�#ҧ�u��sU��8�\��8�D�^C�4��E�r�S5�'���vl�V����`b���y0�t��}%��++w�U��
H����
�\1C��p9x��)�ZRsP��D�7�)\h�r�,~�[K�r��}�"���	? �!蘒���=�/�g�Q�\��װᜣ�)Z��&>��8�uIA1�T���	�}�/Q8��H����"�x�0��m���\Ꮁc-��C�O�t�x@���.,DH�%U?ҫ�H�%��Ԩ�)�����8)�W(7�������&8�C�������'���Y����d��g�@~P��|Q�Xp�`&4�D�c*xe��pָ�U��L�	\:�vV��gK�\1@�������j�����BUI
ܶ4(�!��[s��g��E���c\� k�F����������cڐnT�~eXڪ��w
CM�\�j�ѵ����@J<�A�h*N&M����'�Y&�Ƌ�f��{��fa:IJ.H4��Zh�s�|W�޴��>rF�P��ī��+��30�tq޽�T�ְ�#B���J��^�ЮS~�D�[���!�R�_��76���M AaJe����q
P*�W�Ka=�j�m��\W�x��7�IX�>1���.ɒ�}����Kw���:cqҼ�h���T���9��Z�
G�%� +2��� ����\������d�`�8���gfY��ѝ�ٱ��2�wR"��yF��=����ָz��L�c��5&�ل�3v)�ӯ-��Hp.4�ٻ�+R��G@��:{j��S7�jR��:�	�Mh����uC�UET Y9E7��h�h��n%�:�So����$z�3�B\"���<Q��g�m%�5���ʚ�u���T=��p��4wܸP���ģ{����[�Yb��\���2&>��� ����_-��������ȡ�MU|�9�<��ፔ�x2�>7~ng��i�dIm�& ��}���}�D�[��5B]Wz0�zA���=(��IHܭ�uɠ��-B9T7.���f�ُ�b��"p�][ ��0}@W��*�ZbFӎ���"/���c�[���ܙ�HݣQ��	:_c&���K�偃}��FԫTc?�<3�^�"�ݳ^m�^������Ǳ���T�PK��T��E7���{l�.��[�t2����^�ځ��r�����i�e+_�Pyt���7��~�u��7Pœ	�f	BeO԰@ӗ!�`F��N���*��y`F���MP}mUw���ԋ��Ys�QC�H���A]}C�(��-��2�Dwd�-�z���g�\���Sx쥘���RtA��s�*B��>l��v3�H��2�����K�Mj�#|��лQ�M|��D��%���G��dpHu�Yv�N��[Rrx�>���f�_(� M���Fn��x9-�k5�#��1.�:��d�c�����g���tJ�>Cch`�p�����Sh
�&�J��6�%���,A�:�像������I�j36�a;�%����� Tڊԗ��{
M��B �_�K��y��q�O�_���w�9:PlJ�E���ba��:�q\��u˗F|����C����Z
pVj�~\��ឋ���`s�/}�~�}2�aa`�pW�Eٛ'�E���(��y��1���3
T���}���툰+�y��?��H����1��H'�Adϳ�^ʴ����*!+ �� ��K*9�T�������s�p�AC�m״�.a��
9�7(��]I�� ����7�\@kъ׺��E'&���Y�"�d�m	�dH��O�N9�:�G��5'�Vԧ�	�~H0p-��T�t���i��ʹ>P(�*�1y8A~���AkS� d�<��Am,▌���e�ZQ��o���u�B�]k�sޗ�ᢗ�S�2���=Ķ��Y|=U�?+���8�};�� �����Q۬j��|�]� 2X�0��[�{��|:�Sc3:,�&�-{=A5�.z��A����7JXU���³[jT<* 6��~B�?�m$t��Or��É����Nn��`�~c�����f��U蠔����p"/���%'Al�oh�2�|����VF3�����ӌ�O�<?�!5�!L��kn(D�f!�.�_ɠ拊��s�}x7b�sߋ��330^	�ͱy�qSvJ��D�����#;�6�B�m� (�:��4 O�b�Rы�����A�1����rͺ0�	�"�Ųŵ��k��T�ȵu�}םFF�|�b�2ݝ~x���h�&E����D�d���c�3I�<K�<[� �h�[������b���\�s�<���3��B��]�.�x�#)��_J�0��5���_��Oi�]\;��%9:V�'{ ����p���z�� t�]�xH+�N��O�ค�U�*����m��4�}�|�o�bN�{[i[����r�-��lũ{�V
SZ��&P��,�e�N�Fwܸ��~��,ʉd�['d�'����)8�o���[���uf����b'e����X˼�?�|�АZ�>UQ��;�A�JP�l�&�l��P�l)"N��@o����� �l��[�8P�8G�0�E��2��z�}T^��."�~.��l)(5bn�,�z��4�i��sj�D^�?f8�ҷ)�?;�7��FrrD�g���@��X�CWw��Hc@��/B׎�v�5�n�Y����r]/}{��1B���Oq/o f�*���k� �u���B
i�TDj��?{��Y$��d衮�+�l��2~�������"��:�0�va��F��t����!{�ERT��������x�E��5��ࢳ��К��O��sR�9Ҡ�֘#33��_��%� 8?�V=��Q8ߐ`
���s�SRg.XQ��B����1�>�|�Ă3�=ض2՜G@H��j����g�h �Rk1��2M�L��~�O~�|ȇ��%�G������ ay�%�C��Kﳈ�/E�gv(���[��6t�nA���"-�J-q��׎����	�Rh�.ӆw��N����`���r�<)�8q��~������j;b�1kԈ_r��
�2{�RV��qYC��3�<4�kV�48�a���zᶴ��#A��F��A�GJ[�H�qT/�q�?#(Kszg�
S
�Q�s��r@����L�_$ka��z�<Gp�lt��y�����$rN���6��v���^��T�1���`�{G^U+&$����>TDuRۉ��4	.�eׁ��2���C*�x�~!�o��1҆�cuV�ݕ��G^3f��W��:���dQ����esMk��7$xk�{�'��2�k�X��X��o�.��$/=ѳ(�\֑ ��\\}����6�uo`A���(��0�<�S�����KY�?M$����Xs���u�YZ!J��I�Mr�B9��`�}�/��[<���)����9�<>+��] -�����t����R�DJ�	Bgꘗ�nR/�W��&��JB3,���5r؏�j����
ƒ#��Miò^���%�B:6ɚ��է�Z��W��>�7�Q�W��"����\�s�w�Y���e��n,V���ނ��&�y!��g����Qe�a�aNR����A��5a��Rdj!��O9S���|��>d�x?ڱJ�y��8�=���o_��c%��J� ��#c,���* n�S�U��]�i����7$bD���銛�g�{ȁ+�0���j�c�&�)��~^{�1��2gy���+��;��E�E7��m]��q�o���	�C������}5��x��7[�_iv�R��g;!��V�0�G�E��Rf�[����aw!o@,����#Ȋo���� �SQ_���j;�\ͱ���9��e�ٹ���ݙ�+��W�F�!�����b���g�(�ez��<>��p���8�c����2�I�my���_�I�550�x�W�&*4��6�N�5q��Mv���Of'��Z=�������iS(4�s �q �eث�$�����h�����m��������3�J��h��zB�'�\���%�Rsb/�Ah�n�� m�鎐0��em��@'�Ƴ92�a&I<�Ǯh
�G�Zg�e��C5�e ���ԩ.�j8&IX馚f)�.�<:����<_�@�J}�l2X�R���[lw� ˺9�7�Aq��-t�������g�&�cr�]ć`l�l�*�`�'w�(�΁��k2h��"�xcwc�+8�c�8��|e��P�/*�7�V�߽fQE+�w�-�K����9_���O�^A��ն�*��ܚV{�9 ��ڈ�8�g�O��Ц ���0�)�;N�߾"W�^d#ea>�A7�l<e��c/������ڈ��;�� �Y_���\�Nr٪J����bUr���T����އ���Sh��S�C���9��:Ɩ>AD���G,�����/��VD�epx�8�`�r���1qHXj?S��H]�������IiQ�?�xʑ_��I~���~ѣ�D=��㷻(�����t#�CE��큷�{�i�/Lk����n����x�����<��fCC� S} d4�j��	���3�=T˃[@k�k���"״�c�Y+)��"#a�Pk�4;��vb.υ�+�s��|"�댌|#}��;�"�p�ӳЈ����V[�3ӆ�.'"��ٱ~7m��ʘ` �Ngڏ0^utx�}x����V����{N&�F����WA�+���Sܦ�캏�AʜDn+��65޿"	����$��i!kǜ��Z��O�������ob�
R{�Y���m�!d���8,C�%O��SX�M�J�>K-D�2R@C�+eŉ@i�Tm�sZ)kD�v<p�6�Pv��Fs����ū�!�i�0��~
�qBw��˩��N)��4�lrdTݗ�yPt拝��q!��^��v��Z��^�K�ϩz�XF��DȪ�c�`777�
�6��83x�]��l����@j����������8��M�Uf1,���Z��Y'9l/n�~x�\�y%$j�����3�O�V����H���4�J9:�H�j��vQ����צ���R�ǧ���R�w*j�W\�f����͙�}5�p��x�iR��KcC2?�s���Ϯ��@4�g֥#�%�:uX�qwX�	��}?�x��!���lJ7H�_"vhe^�#g�cjn ��>^F�a��M�OR���1[ʳ��h�h=�k�V�45����˽R=fG��@g��4u������u�I�kX���L+�p�ē��&�>�NW�����������Z��i"=��}*9�wB���#O"�����F��eųw_��(S��9wW�-�u��$��gE���c'��k�{��m�L�=���k���&��u�'8m\�����d���*�Z�?�_���ߞ����
��;� �\l��&���-O�hdB�pRU��TI]`�:�	_�b�������:���n}�A��j���+}*F�^��[���Fy��V�����õ�C
!���g9����+�ei;�z;����g8���W����YiDV�)�� A<�^i��A��~b'u�B8 '�xsrq�9�!�T*T��L�|~�s�*
A"���J��|o��� �M!�&�l�WF�~&q��I����龅�06����A�n�AO�4��
wi'�ˏ�)��`<��~��6yΦ�l|v�ȳ���ƪpN	�TQ�A�E��F���Ny�$zR�#X�~��w��}�w&�f��ߋ9m���<?0M%�#�)��*�)�r�R�-���I'�=+G1�`�U����� ����[~J�N�9<��6q�N7�s �����dYhF+5���P-���p�fN�-��2��m��@�k�9t= �՚1<�Z�
l�|�]��Ny�z����yDt�M$�z�T�]%7Z�Ih�y��q�p���#%�Ob�w]u&�ņ��܀�ll1��`�K 2��r��%�h ��:<�����l�5�dk
��D� ���j��~N���'V'�zan��y�ʂ� *N�GY��T!U��UPQG�=�H9�X"���5�[�9�w2C@R���)u�$� NLW��o�<�.���v���q�ԃl�=�/Bj�t�^e� ��mg�KBt0�?�Mz��c	N<&;�M����.K���,K���gg87d��l-��A��k$�ц^�MMPE1)��KE��'���D�OL��V�p���9��8��k������7�a��r�U���7=�d���g�v��E�UG���-	x����QY�R	��r9<(il{{�8:�E-c-qi���,#�a���Q�I��9�ah���-".�,j�"4��Y���P�f$ǰ�&:bה�sC�SD��df��fNy�bE���IM�vPMl�K[��׶-;�.��${�R�m�;���皃��?�_� ?Q�����8/� �����*	d�&�[�?gP��r#,0a�#/G�m�t'��ߏ�} Y���0�RM$��f�O}]7�1iM)�������,���w�l�̽�c�gb#:�4At��'�v�K�Vo<��?���wO�7#��3&��#g;�A;���	�J�ο^���;y�z�u���Y݋��k����j�G.y7U�N+a����_A"Zu��v��|-em�}��
�� ���a�ʺ�2ǲ�b�ѯR�lTG������x��4�[��q���R8P���a�(e�N��|)�o��0GtsB �uz��C�Ug�#�}�	��ե�g�XS�����;-��K��������%�⊟,gwȔ��Ũ~%���k-�8z=�\�[��.pR��B�0jl���8�K��D�!h="�>e<}��u-ё���l����I�-Bb��2f%�[R�(L,�+��H��$�^��vK"q��ےR�rU։K�m��q�e�樫� ����b�.�l�*soJ�4 �9�� �$	Bomf��.�
l@��w_�4
.�,�;w�=���<ƕ�0��|:�x�	4����,�H�Qx�~;e8��͈���ֿ��sa��.�su*���|vq{�4_H��8�%��2Z���
���q��A��p��{&),V�|�ZE���aD�q]4/J��j����ˋ�}����œ1K��he5�P���!�A2����P���n���h�I����st�?��T�,cr3����Mp=]��d3���9t��i�&�y����>���-�	�
����̥	���Y�X�.�E��z��,~���J��9e�Bv��V�QZ~�Y�YQ��"������ߋ��a��')��u�����J��V��d�fVG���y&�k�_��;J�̚U��쪦Ѹh�k�8-��Oy��z�w��O��tݫSDd	aN��[�}�%�_��< u1~��}�dV�f9�R�Ӆ�`�˦�ߔ8�nP��6u�|��A#�c:.~Aai��*j�y�^���IeZ/@3�Z���NMd�Z��|,%Ն�����z�ֺC2�c|8�1?������*g ����Ż�n�����lG�A��&/g(a�Q20 �< $�}�����|@�YO��S�:�~ѥ%�^���v;4�O!�h@�.ٔ�F��6��Q���,ڊy-AD;��ʰ�}'Ig�F9#�?-��*_���)�{T�Ω� �T�+�|�w��N`�ܯƤ���9a�ɲ��7M	��5���i澻�$�
[X�Һ�S��Z���*c�X�CĹj0�%���4���h_}�� .�դ����2�o��=S�ST�]¦ � ��>,,"����U����$��N`�E��Ԯ[�0�2���V�Po�;���R�<� �ze�[�ט�23��t�?ـ���G����#'=��r*<6�FBX{=�,vh�S��0���z) �2�G���x7�Tͣ��J��X��B: a u*�4�Qb�-��j�g4������-;��| ���e2E�z�9Р�S� �o>�YH��^��~ʂ3*�r��Mͅ������5=��<�@��_���Z��Gg	3�5�9Z�{z�W��	����ʞ��B�2�EYtO�g�Mޘ>?Kd��AK!��fE�m͂ݨN��u4������^�t�C�6�R9]����/�c��R��1�}����E���b����j="�cM�Z/��UT���ň�Ѐ�j�;�;"��`��7�����`� 5�A� a��I�$�HDzoH݂~���J��j1B*������.'���{z�V9�����̽⓳f
�In���J���fװ�r�������ݝ�M��=|D~XvϮL�)XR���1�*ٺ'�z������1({y�i+�Z�r��й�{aB�ju�̧�M���<�}Ȣy�u���R��R�>>�Z�jQ!��;}�ݧ�H�[ � ��Ŭx�@�r����/3ٝ�@8�$v�t�j�ꅓ�z[�w鹩+����T-�A^����[�݈N�V�}�^�h�d[�h9�1�����w(��S C��߫k����_�S��c�Ъ�w|�
�=�O&Z`3T�A�C��;��	��~�����i���T�,r�T�-�-��ϒ�^���E֎n�&����͇�}�P��4�w^� ��!�e�jb��2����=$
��O�u��F��&%�H�&d�,�Qa��o�W[tb�(�Ą1_�o���[k�_�x�5{Y�4�N�}� �h��5{/y (�����)�ڝ�EhC<F��e�Ƃ�d �l�^s��[��.��Ţ���M7���kA�=p}4q�}�[��x|��W�`*��V�"-p,�4��y=	w�\^eX;��^P=�ɴa/o��vMP�m*
��E���ߓc~�uV�<��ĳ�
���t���(�5����ܞ6hJܣܴH�%Z����@�V����ٺ�9����n�L��"[���Uv�䊩bC��;�q���vq�D?��+��]��������pO�(d��,e���^�d�i���S �x��!��N����~���{_�����ߥ�R�ё��������*��KQb�,Nvw�ZD�Wq�4R��	��tK�B5�G���qqZT@��1��sd0�Mݘx]qz�Gg{�����)��ަͱ=5���[RЎ�B	���n��~JQ>d7�����tD8�fqϾ�M Q�p�[�0Ѣ�����(�U�rԅ�B��4Nw�Y�E9C�0V������4�{�z���c�m7~%@�'����y'�G�I���F��DK[Ʒ��h�c*|hx��+g$��R7W�\V����K�z�S�H� �`�6o�FG֮oM�N�%��rŧ������!�w[���*㴟V��Q�/T��*a�ـ_�rH� ���pm��ǟ�s\��D�8���ס�3���n|�!v
�Փq�|�U1[n5���%���YM��0�1�ȧ��+��v�� �%���Ou�|D#)d�	c5$yy���^��
<yV��/҉;-����ecL�5���հR�F�\��Dd��X�'���{dMI�2�]_�W �:T�`����T4�-&�x����s;��.���T�%�c�	�*ߜ�P]��J��#��ǃj�n�A���fS�u��"�.4a��v� ���ē.)��8�^Ґ(�R�㸚��*skM�G�F�S�L"����7�n
힉.J�i7�8\3�9J�nz�
Ý�7��F� ",��'�@�S��i�O����O~ZtF�]^���M��b3fk���{J$��=+G+�����UC�H碽�ev�y�
&��+DD�B�5&P=-��N���x�~���ة��H{�`8��*V���m��B=���2X�� -_��!�� ,D%+/���OU2����1�?}n� +�5����N�G�	ur�C��$g�@�ĲwV�:�qO�M��Ҿ��yh�5��x"�%�xI-���7k�3�l��8ˢ��[�/&$~]h�� QϽ{��Ff�ΑE�kg��0�yaå�0�#�d$��l��2�r~�1%�a�y�Ud=�������KY�#?�I��ߵ�&�]��nD�l�@�&Ǘ	(}<G�qK��-�+I~n�K!ѳ��v(�P�#K���&�f�N�r�|�}�k��Tw�Lt�)�[��MnlX�r￿4�R}��&u�Z؂�WMa��dK�|g[,^PU�2kI���w��V���5Ey� ��rZ#�3/���c��'��KXz2��P��s��,�,d�X&�o��8����<��!
h`��m����T����'���֛�4�e�����,����3&��}���`�r8�c�moo�4�~2L��0I.�,[��a_���܏\�K�눼� u�~v��G*�Z�:Ic�Q��=�ƭ�������U,�Z�H�,{Sὄ^�ix�<7v���1K��Z�Ql�	�^�$ԝ%m�e���YK�`Iߗ-xh`��=�B�I�[�{�@����u3e��C<-p�9���KB��8*���ׯ �y�m@��k��Ur�`%� w(n����+�͚���A �H��aPXbԞ�ތ[%W�����
hj��%,U:��d1G�c�x��74fJ�׆DDs1^�MW�r�߉|�A����ED���L��Z�Qq�3R�&:.&��c���ϲ�-G��B)�Zʩcٷ���݉��q�֞����9��%{�L%��FQ�.ծ���]�u��c�5�lL#��+��J��ɢ�&�r	��Y�R��d��%p�$x�S��2x]���w'�\�i�UV&&�(���3m^9꒪���OIdp��J�KF�;�WlSR:�O-�\�P0Q�����<R͙�m*��m���Y�`�sתV�=a�;g��Pcg��)���ň&���ӓD�:G�b&��ਙ��,)'��-Yuά����������W&���c<�1Zf.��k8��{�ô�gu��{4�JV]�rM`���q1:}V��KE�ϋ���i����V�tY�����sn'���������51�����M&"ޡ �V�<�9�B�GLux�U�"�%уT0��t�N4a��Z��|lt3ּ<1ұ��1:�ǽ�q�o�2dgA}EC�� a���a����|/=rj��pi3��c՗e����5`7�y�i%Ճ�Of�F	�\�Q㬵or��F�6�s������g�ᛄ���Ӵ̀��
�+Ye:$���57;T��c��?\��y�3��jUک_��ȥ徙��-{9�M�,f�*]���\�	��騢!~�'� ��t|C�:��	l�S
�&��h����yh����9��L��o��߀D��q:I���QD�I�ӭ�E�e6�Am��3@�/�b�<d��=���S��R�x
�������PxLD71#�����8n,ȟ�5����#e,��#�P�i!A�YoP�<��OAԦG��+�x��gZA�+8�C��.�肞N����ވ�z��s�M�<����Z�!�$9��g��_�/t�X��Y�Qx�A��k+�	\L��!�q����7ʖ�woq��r�z��F���.�b'�K�FdeP	���8���
�|j!IQI�Mw� �ܓ��6�k
�+XO�+���;-)\!Ōp5'Y˯��=���N��k���7�������uh����h@lI��B'�1������x =JP	�œ�y�Nb�I�$P��������)�|�D���8Z_�ܥc��)��U�6]������[���@Q����T�-)n4�^D�4�����R؇#���]�HR~���{�vʌu�c�&���F��ڥ'��K���B�6�rI(���޺K�-�,�p��i���J�̷P�oQb"��^�v�b�E"��j�'e"m%Y:�y�6�W�Q���]xY�ydÍzq��p] %E=�v'�/�=gK�ax�,fXKe��<y2f����cg�ó�A@��@SL���Q��¯I��vJ��
�� �L�ʪޟ,+��i"t� �(/�v~��V&���^(-��p�`%�#iE�d����g�l�,Q��\��d��R�\�鹐�@�gL�}$K���bU�)�4�9h[i��%3���H��Wڜ6��s���OA��K��}�4������g����gC�1Fh���𶔢�L��%`u[V	\��� ���[�F�c��::���_� �f>�+�sS���s!8���ցx,>n_~�xɰǟ���������RG�Ҍ��b���!�." ٪grh�q�:Sp��1�U��v��W�jOt}�br���Fs��Bɳ�iv��4���ٕ���ڽF!��}��+W���ϰB(��f��u��'C!��/&_E:I��� ߶)4��k��[|�e�+Ə������9�^i-� ����.I���+����۱7�=m����VZ<M��3
�+�.�{�V(1U��N��m�\�ꏒ�T���zv�`z���������Q�uT�I��2���YK<s'M��L8\>�E����P[�]1����`2�*�N�MW�
K��	��'<+y��P�F��T��V�I�|\m<5c(�X��y�,!�"�9�Y��^[�(���91x��>i�*S�����u��D���!�xV�#�a��L��s��ؓ�St�V·��F�Z����vlcy�!ݮO,��h��I�uI��,R�t�y�QR[��"[���Y���SĤ��L��.����[���`)�5�=�h:�^\�
�W.#�ۼ�b�޺D������i�����X�߽h��Yv��u���]WUU�q��Kt@a1�e���J�&�k�tY(�� X��H��� �f��D��д��!-mxܔq{�u�堈�>�x�Q�	���p�X�'���	J���&�C�X�Qn&;�~�d���z�x+KevhtAw�n�3t5X��e���bjh��Ϝ�a�� ��p�^��u�B^T᜻*������s+���Y��x��+�o�Gr0>zm�sN������b䉹�����(`��f����wA�^d�e��L�fV|I���o+g��?E�'뇥�l��޴�=N-��^<��B귘�N��y]��߬ξ%�#rp;�nJ��@�H6�}�nj��en�UYp8������%J8Y����֍��i�5�Ḝ�0�ysP�<��ϳ�pXt���)���P���]%�����N�#;״w"l��Ü�Do�͕�-�>����&��x��@����v��0~� c^����>�h�~���/'�2���so���P�����%�
��Fqԏh!W<��d���3��z�n�!z�#98����T��@��[t�`�a!�jM�)]S���WrS�-&�\; 
�����]�l���T����f�ҙ���ac�O&�.�n�����*�%[!N��f<%[�Jx�ɇ��]��R����7ԙ蟍j�z��
��Am��͒%uT�<�=�Z;p�(�~�*��&�v�Y!B��#�{��18��By���&�� [YÛ6��F��3цn�i[� �X�uc��S�����x%'�]US�����r���X%KqA�	�$/���"�l>:���D2���]�T���ldL�Tc�����r�{�}R-�F���=BuQ6ς:'�1����*Z��e�/!QCs���Y�������S_i<��G届��i���	R��`�(�'�E/�8���V?_�&Q&F�	R�z���n������hԜ0-K⅐G�����Z�5������_wAH`;a�-�TL`�~�ǈ�W��ױ:��042ZJX�'~x���BZ ��&hު5*������W�-w���I�Wl�|�i�A�x:��ɿ�����!歚o�R�"�J[��E���yE��'�!������f��{�Q�����Ϲ�-������ ��z�<|ySR�B]�ͧ���EfhL:��N���Q�_n;������٧#ڲ��O�1G�7�U#��Jħ����	׀�e�ڶ��Ue��73$-:#g%\8��%���3}�>@5���֨x3ܓ�t���NTE��e�hdp���z�UG�֎&��m�b�^v���8�}�o��6�����CP��<�'�ت�I��2ͺ�yv�w���t����IjײB՞	o�~ި�Y3_S���ڰ~��N�h�d�9�L;��ܟ
��w�^ɣ�%)�F[y��0�q\���}�\5�g���3�n���[��	����kEUX\k]B���#ࠋ��u�ԃ��xlϋ��!�Ⱥ�@y�_ SW�fO���Gِ
��7������.�uԥ�C���)grk8v����d��uU�Vޯ[�Px[� F�@hkY������ �t5;�a���V �b�=��<��`JnD.�ݔ�"f���>���̰�޴Wٷ���Y��@ ��쩿���,�%����9�jȶ�	�sĂ*�cq�׉���q�L�i.W�y�K�;����r�'U6f042�7�Yi�h��zɖ6yc�C�:�kG�\���8��5r�uH�m~�4]�y�65��䏧R:F�	�Ə�*�v	��9�]xJNu�栜��ן=,X\���ɺBu��߶�1�(�$��zC<J�%���G^�Ƭ����I�|i���׷��_­.��Q�����
>K_&�r���zi�H�C�\�"C@t�&P�(��_p8�(;��=��G���L�L 9|JLO8����=�J���[$���w��$�5y�r�S&y|����H��qR
]Q	�!1��o��3�����mf�D�On���H��Ȥ<���l�u^EHؑ<���W�~b�Ǳ�(
�S##��i��~���w��J��"jΥ�?��*��
�X���'3����#�,�}���1U����m�w�����0u�J:�b�-)[���bq��}�Wխ�sܘ�̤�@Z�a�H�2',/�0&�r+�q�e1���%k̈l;D֋����ty<F�NJ�h.M6MB�"��l^�^�Җr�Nf�ag6�~�WB:8�T$�F�n㹞�O$l�\����9O6ЬC��D�w/�P�K�4|�. �2�W�}���c@T�3��Ta�p�ж#q�G���ٵ�`�3 <C_���@&������6m�B����~���e�� ����g*���ԭ$@���619i��>�b�!S���vS�RD���?.�z>�}t1����h��ֶ�m.��T5��w��0�V!��i�J)�tR��FF�-Otȗ?�KϱD���8�K�o���}W��V��vF�U���W�̅�R�MnÒ�
�����2ї��?��H���Ϭ ȫ*
�����E��a�_#�rנY�4_A/�i�.`+�ۯg�%f�j�ۉ����{aN��p���������QbF�a�;�0+g�!
�f�+�qa�Q���s+��^���ٝ����AZ���SqrN $���Һ��(���Y���5>�B�_�V�qq;�]�@3d�����2v�cN���i�_��`�`�������`�>= �V�����d�'Pq�'�tī7\u��R?	�H>���+�=m�>���V�I����5�};$T��5�ۈ�l�x�1{����cXxr���R=� �\?	L��%�Rp��Guਸ਼���JE��qw`h��Z4��PK��$�	y� �8���1�z%�R��1���T�����yV�V��:!\���(�;h)8`YD��$f����n����y�`�?d�Lckɚ��H\�w�:�v�U��Ze3o���J�&3J!�V�G�Ϯ���Z��8�}��(�
_���@��&�ܩ�-��|(K�L��oB��\�`����;��-܃sk�.P_���yҳH��:�"g�)�(�B;��uS0q���\���ʠw�@ �͒�E�,N����x�g�_"��/��>3
��z<�����C��!�`v-�Tq����\^c��U͍�*Ġ�ւ��d�4DhZD���M�ֽ��{�pIR���ӎ"��
�1��_v�$/�2���kQq��Z�8H]F!��Y�7��
0^:N���P��A�R�k����D�3�C {�.Y4��3WO��ͦ7�\��b�)�.��ix��%�*�]p�z'�	[G��!�����=���ݧ'��K.U:�p�Z�5&d���f����5ef�ژ9��;�a-yq⮲�d�?���O��T�~�����Z�r+U(�����ؕ��%u�rM�	�s$$�v�=���_�n�U&���lP�~x���9U,îx������ ��ʊ�`Gt����qx3�}$��T��d:ʘ{׮Wg��i��������?T�1o�i�� ���) %M��b�tݠ�1 Ҿ)wp�����u�Dg��$lnc����D�͜Z��ڴR�6��QJ�y�� ����A���}�O�c��:��(���� �Y��q��������Ooj�WFb��|��'���	)�`�\TE�b�=}����n��X��9==�#������ 8��~.�@J�Y�9�Q�{��-FЧ���"�����cĪr~�˪!(B����o�U����iO�n挃�*C�������T�$>�������E���u��Bwvh�5ë���R��]�̌e�Qμ�f/�[�jܗ0�@SNc�h����~ஓ\@ �3B�/V/jp��9�g/���~$6�d��|��Z �]wBz��4��51`� E�y��</��
-�<Q8���qJ�y��ӥ��V�̪�A��)bn����\�H0��K�=�g�q$2.�8c���4\V���ō5�sf���w�Z�;Kn��iᙾ�&���,��,=�~c��kWW$�|�#(Mv!�hvU;
,";R«��\��\��������F<ᙋY�@�7�c���
l�d&��a�x����NC+��mߟ�>vF��Vf!A:U+�_:@�=�[�{�L#�=�\�Z��܂v�ȼD��X#$ަ���TVڭ�d>=m�s�;vKJ�qЩ.,^�&k��t�⥪�ƃ��Z�T�-�F�4h����b��S��%:%
C�\ ��\�6�x�&���3֞�w۝�t��8f<E�������PҊ��^B7v���+͙4|<2����Q1[�,ɑE�<��[	�?+
Ww��c��61f�5�N�*F.�͗t��o��c�K+�- ���oq�D�<�^Όn���b��)�^�6��+G��a��HQ6�Q�h�kޠp\#�~g6) ]?�	64+'0��E�_�Sg�a'i�5��Ԉ� ���Y2V/�$������,8��Xb�9D�P���JR�5��\ �7y��K��|��3�Q�����/�V�v&}���w�ǳ���@m!(�g~�_HlLglZ���(ț��#<�Ѡ�N�ߧ�	'z��Jb�1��!�R��P�ë��o���9�!�5pPd�'�L�ҰK�Wr�H��o������>��3���.��,�.5��?�c\���p"�ح��n���h����-r��ڷ1��Kǉ��`0w~q �zo�[��(���O��)�.�93Oc�/Ot����-��e�H'�[�~�i&�4�7g��F!y��'�e��x�:�I7�N*�@8���x�5Ֆ�g�J�1]�7�'dK���Qsj���&β_.]��3������3w1�M|�+�1(�j��Y#W�5��u�R�-��f�YR����~����
��j	��S|Q�,k�˜�������%��{����5�\m\52�v��Z�V�=�b	�ؘ�5����7'�4���O��W���p������D�qd1��U�%�R+��?����K[�����ʙBTf_A�ë���o[o�,����{p*�]AB�>��͜��ƹ-�$�st�4�\����<��s|�c݄+�`Խ7����B5�WL��`2p�6�JܧZ�xAK�<R��3��8��>݂�����np�!ܸ�د���+)^V%z9�!"��{�����8Y���G3͜mg	YD3R�֙qK��Ǔ�R�  v�"���e��<_i��q�)/o�3�O�Q��\IP���F����F��:��i*�>M6Ι53s%��,'3:%u���Mȷ����.X�S���� ��]����� x�ޞ�.d s�4��\G
x`��n���<xXa�8��2��4� t�Փ���F�,�-I����h�����8��.�sx$.8
;7�:�JM�a,ԅ�_�T���=��;Ö]yo��9�4�.|RY�K�.Կ���ح�bL*�^��^O�Gw���B������zd��a�3&��}v�D��$-��:u�"(���ͱG��P����@�Հ)et4*����ݷHvmڼ(�vu��$+P��x��G;O�4�C��߸rY����P����1���O�2�w�zj�dť#'6�����C�[RY��*;2���ukP��*Jp:0��nV8�V�Qi���3���.D`�"�<}0�\����i({�PE�C�{v��q�%ؐ)Q��Q�['qͺ�"
��#�/�8�Rjxλ���4���<r�S7�g}��3��ڮ44�o$�e839ѽ���2r�ͣs��'��Yˡ�4G��Pݝ�*W�F틡�]h�y�4�0a�Z�ݮ�~H٠0��U�s7�Ҟ�Zq�C�P�^*SL�V��(�TC]ǣ�S�-xR?��f ���B�t�x�Q��h�j]���ݗ�C��|�\(Ҡ�sM�R1ԍ��ɵ����'��zKJ�A����vF��A7�U�pr����7X:Kxᑜ�b'q�G͢$S��Yn1��s�桉p蹭X���B��lӧ�mi�}F1��%�UCԻ�P�h���i�foW����۱Z{�{a����bu_��˟��K�GA
V�S����kR���~qX�(�E������܈P���Ekd����mJ���������7<�����e�ڨ]�YsG��>_��0}�G��oj���%k����v�����#P#��߇S����oX��ě��������m#���t́�\�1F��+Q�
I���'w�؜KIs,�d�ӌ��3�b�lx��q�Y����º�K��dpZ�F����+}��"5�a��߿9��+d�Q���j{�\R�[�d2��X��#�����4�b?_�@C��������է�_^p��Җ�m�Z2M}ΉNP0T�7y����vV�����)�|�s�jA�H�������@4�;���|�n�J~<N����X'�p��lf�|X��BE��m&��c���-�6P'�
�K��Ԉm՚>qN�����bg���^�������L`t�ɵ��V���/{� �\�wȢƨ&~I�U�1� g'�?��B�4�$�(z�����pf�0�)Ϡ�:���+$�~����4E��q���_��X2���D�ep�XN�obb��4��x�@s��?P0�ۖM�/ATfD�]��� e�u-le|�}��K �U0�e�:?��%��kfԗi�{��`�cr�� PT�LG)�QD�8�7t�f��n��|Ut���XZ�Kϊ�����M�s�f0�w�9 ٲ����/�o
����M����K����Qt�OV";,��gx;xw�[�9��S̃��ײzt���~�����|��ZE@8q	�D��n��>S}V9������/�9�>�s(p-��3$�n��Pt�<,�7���4f>$f�~�m���&�p��� �.���;��o✟)N�i��ind~f��p���sBbr���fFU�҂��ځ~�3;q�#۵��ǧ��G� -����J�pk��Yj�9�����&D+x�]��8^�	!!������*���������nK%2�@�zQ�K3��K�$��J�������e�)d���/�	�+�9���C��'O�Ηm0��[�a�p�x���8��=���/���cLO�:'�Ltc������}��x���f؞
¨L��Npͮ�"G�cO�E���J̟nI~�6^˛ ��6O�1b=�܁�C]�;]bV�����4R�Nr*��P�H\
ڱ%��v�>}Ϗ��`�l8� ��.�~�����G���i�_�OR��Lz,�l.�S����@Le�%M�Mޯ�)xZ3xBw �Ù����qx]'ѳdۛ�S�.�E�0
D���+�Taqy���B�v�f��*�8/��Q�:d[?���\/��U"ʀ'���[�)�u�J�W�LzF,B�!��E�0��e�A:��O�}Y+�����s��Z� ��*��D.LI�[�.��-�zn�A����7��^��F������mjK�ǵ!�f��D�ku4Q٩�@7Q9�>�P��iZ�ʂZ�s�	Д�O����nc����S�7H�dJ0}N��$䗒�VX��0�D-'��3��Zk�<�\pE�<SdĹI@�N�?9�|u�c�X�%��>�ǻEf��L����J���>�OlѾ��Ӵ^�{��ZT��[k������w�Z��[=߹,��$�u�_�|������{1.+)���@,�Q<Շː�mW�D�i*WtG#=O�5�.�B�*থ� �Tm$���-=e��L)�%���6th�AO�|k�{�CASvO=��c�o7���-�@�}Z�W�yj|�-a�
l�
ĺI5(T�!�Kx�D'��45?0$Iq�`�jtFp_��ZR�2�C�Y�Es��o|.p�.�n���Qk\\脅{�#?��E24Z���o��9E$�>-��N{�Y��� ��m-�sϕ�V�Ta֚儊l�t��CU���Sb�s��MG7�#��8��'qc���T{�W8�M0�
������h���ta�D������y ��П%�bzE��羴P�X����s���3���Cu�\Xg&x7������XUkS�R(Yg����Y��U9�qWT�7/�4�]�/A]�S�r<�8�#9��f��H�G���36����,d�"D]��p6�8��j���4{��y�ܳZ��4���,�P:$S��~W�!��/}l�(}�P4+���JV'�8���s=��xb+t՞�����)� y� �M�啒'��ޥ�W��O�{w�/�gOlm�µ��q��:���a����o]l=!�ΞV��|�Ү��b��)Ka��]�7�@��_ӝ"،�'���0�{���*�q/6��%ۦh"ʹk��jreM�2������,
^���c)������_��>��?�^>�.�+�;�\��+�^�7Q��&t�Vӱ3l6h���W�u���:��EԨO�qt�1�u�F��ۗ��OA-iW����|���0��hi��;��RTU5��4<�>
Pȃ|(�Z�ލy�3_ׂ������P'\�Z��+׿[H�s�]��� Q}7���ɋ	�E�w��Cc1���k�*�.�-egGc"L���w�DqX����I
�.�]���pFSÙ�=�?�6�)N������]A!��u7Z��C�*�n8�<��kÚ�2�K����Z���Ѝ��#޳��6�L((f�;3��[P�8�1��K����7��JqLb:��x4���u�'9=������>DF�U]�"v�^�Q�>�Muo�x���܊�ڰ�'��E��m���Rh.����O�D/�eɘ1
S���y�x 9w X�Zu��:��
����uJ�|��l3,�I�vò�P�`L�_�5_Ai���+�n���J.;I��[-�r����x�E9QN��4��z3q /8S�� TR����x����c�YCS/�Rn�I�:2��ԧ��R/�]L#�S��&�~7�W�v��\�(	p���ρ�K��V�B)|q�o�Q�]D��F�7?!�<|=�j��L�{0��m��Bnf*�b�T�-|�k��u>N$��3�ֻ|�-V�=�+��J���[���z�	<P��?�g����~�����6��tp3B�%\�Fc/?K|�3�<Q�)$�yO�$�B
$Q�b�&���q}�̔AH�P�1ec�j�f�3h \����
�'��=j��NN|yb���&��B�@_��zJ}�/�T�Jh������<� ��ۋ�-�kg�◘�ܣ�6P?�)�dπ+6Y��2v�2�=l�V���������G��a�3%�X��m�R˨���A���<�m�gm���H�����ֶ�M)ݺ��ծƭo14f䦊����r~1h�`ۛ�?�߅�I�]3s��w�[����{FX;����Y���&��^�C.;�!�?���c��)c�]���|�(d�n#��<*�|`��H�������r�k�d%��0yp�0�h�����o[�O�vw��I����G�0Ґ�;J��:M��FoQ�����6��v�}!�o���{�	:!z�� ��/jDo����Cr~��:�n��@�5��{��&��B����TQգ���}#�n�(���	���W���3V��؏[���j=�G����Z���nr��.o�9�^/P�`���"u��[��x��JO�ɸ*O�2><�|���OO�z��3��=;�^����qږ��1��_�O�8Ϋ�V��3�Py-��^ ��s(*+�WV� �x| Q� �a#���Q��1Hloo����#՝U��'����4$���e֜9����[�2�Ԋ��Ԝu?�j�(q�o�̣�X�����8��	;U��H�w�adtc��lV�qU�5��A�'����o��N|��XiH�2�v�-Fg�??�<���e�~d����1��4�!���$"ps[RA�a�.{�����x�y�dP�g�,rt�r˛�*�W�)$1Z+�-f=�V�@�����~wJxf��Xǈ�cq�6��6�2���n���a�A2/�`�-sX�� �(�J�C/20�\�� ����O�͐���ͅ�m�=8-�U�*�H���h麊>��Ƿ��L���˨�G��QIt�rI�\���QО^��^���JIwI�����A��O�Y0���aڋN�� 
hL��F��ȝ~H{c�)���])й+[ �Մ���3�3�(�#�?�+@��E��ܒ�<F9̚�۰�$���Fή̮��!q�9����+o���{5ֱ�p�N�@�X#�Z�)kF�1��A"^��2X�+拉\���M����}3�<Lr��~���,�h�� �YH <�� �彊::C�_�'���ꂦ���L+��g�LL�`���_����8�>B���d��4���u.���:;YZ��P�¼�s��)u�II"|mK�$�gzy��B�U�~QdV������ںY%�$?؎��O�+����78�̚��&�I��]�U��o�MV:�$�B/��9I�j~,��Z�#�f�&�L!�dY֊�z������ʲ�Y��vȼ�I��z
3y��_�ryz�!��'�D��o���nj���m�-}Ԇ]U��v",�No��\/	�/i��N#'��������b���m��L�{��E �Rӄ }w�殃"���c!���>����+Ӛ�")�Է��v�5�2�����l�9�%�㌙0���D�d?���;]SI����F$��Gb�=��+k�eNq����ǒ�m�T��}�c��t�)�LZ"�Ɗ���m�@��zճ��@]�և+ug���q`9C���%.֌��߀'!�^�������0�b������BQK 4�	�(T�����2KU����V0�z�R��v�YO[	0U	#�<�q9��$<d�?���62��c�oP��11��
����W���4f��*�n���
�(�͙ҸxLzOq��L7�~q�	�vB/j��T��[����-��S0��3�����,l�xw�n�qsz�K�����8��QگW6s�DЧN=����u�G�d��2ڝy���mC��dsi ��F��I�y���+�e^��x�d:�� 3��c�ˇ��'nyL,w�)p"hcɫ�P<��s�p\x81��V]Q[�����'��0'�����u�8����y$�WJ����L����tX��v��c�,���x��*�Q؎��<��ɐp�<�_E���	s�ʒzc�z����<�j<��CO��R#�,]}|�.|��KP�����f���-�K�F <���_�<!ci���"	�?�����MI �PX��-��ʉ5_����}�.$i�#�zVY»8�L�m˲P%S��,j�\4JҀ`���u��u���88���C��eM���N��7�x>7���Uxѳ}�J/�����?��-^�0k�2)��2�.�I���� a��A�30�:���Jka�l�h��������a���6��m"�z��*��_j�����N����
H> A@+dhi�2�ȪS����/V�Ą��'UI�q	fͬ���qc�V����V����⃏����ۍֶ��t'�S)7Pk+�I���U/�!
�X-�%:�M�.��Sp�6��[�="���I�?��ДT���~;	��io���E[xu7	e��\0��L�+9q�g�쥸}���Y��^�H̊�!��;'��_��w{4�v+���A���PJ+ ��Z����x�^�pGn�d��8��=�tD�'��	F�����hf���CY���u�m�{փ �S��E�ܜOu��}cYL2�q��#����hs[�ܾZ�D+t�r�v�w���crt��1V������Ez��0>�q�.���%�X���(|%V�8��$S|�\`�=�	�`�~��]]�H�����=me[� ��D�h�N����ËxO6m�R1��L��CEs	���[�G��NAl	�
�1nܨ���)������&S�I�65�l���rB�U�%r��I����B�3���Od,����g~���|���5��CA�8�^]��[/'���:�d���|[��!�'LKx竦F��vm�%a[V��p\�Ȇ�ќ����'D�jG>!҆u�����-���[��}$���'�UюG�!I
|�Ͱ�F�Z��o��L��s����aP��:��a�8�[����U5�:�W�ѓ�7|�z��S���w7�q��@�,^K���8�<B��*�Y�a��h�.���3�!�]s�T��J��Ք�Y����'�s�$����SU��Z�,�o�X<���2Y�����{F�|�J��J�{�] �6B��F�MN#�Öc�C4�!�y���\7�@O���ͱ2HmJ;��U8��_6en��#�;ۑ�_n�@/<�x�1��>ߖ��&ή��<���=�F�h���]o�+�5=�h��0e��h~ȱ�5�rf�hƒd��w_Pi� !R�x*;Z2�)�%]ʎG��2e@~怦�|K	����"V�!��Hv<��'�v<���5��1�LD�+�˟�/`��GN��!�ɼ����H
s@�9so��X@
�X@�l�e�%�{~k\��TH~|���c��(���y.pJ��:����̪��P�v��rx,͎x,mk���NGߜ�Z�9o��7>7_!�Le;&&wUG=��s��Us��-�����^�S�D�����H"̙�1}C65�%2"c�e��>��,�^%��{��\O�,ϙ�%-i1?��ƪ���>���l��sޏ2z���IQ��b�m9�޿Fu>Ou�i���b${�+���\��lG��i�J:V��$E�y���y�4*�f�m#���E�U�g�}��n�AĂ���rխ%�F��7�J��z�iRݭ�y�����iBʔ�]���3�ϕ�1;�aS���Ocس�]��}9���-��� ����*!>D�_�ѳw{*{��Ի�n�,�3�6=,�0��(~��1	?Z�$���]fKE��{��~�?������LU���yt������^by>�Ϩf"2�J��?Z��1�%%y����q��K�~Nף朗	̜�TW��#��~���ً��Ԍ �YJ6
�fqO��M?s�0uh��o<��U8�'�Ъ�\��9���%T�A�}nK��o���g�ů��7���*�0�����陁r�� $U��D��+�h8�(<�Q:h��@c���e+\��'�����s�?��X] 	1������c�+QV��d�+�ۃ�҄��� ��;-C�Z���Ҧ=�M�b��x���/���[���^�\>�]%֤2�H�qüJ>IvE��ӑ!qFږ��r�	u���W��D�M�͈�w`��cdp�.��X�`���v�d ���ˌ�����ȁ�SMHi�3A�	����R��m#��S�wHfM�+jѽꛍv���tg;B�{���Q�r�#����k�2F�y�wHm)@��qꤘ=�j�y>���Ui�iZp)�YiS���w0�M`\
H���7r_8�]�� ���������ig�\����Bl ��m$�"Tw�Zϕّ;X��x]���p�Q�^'Z�V?�S�|���e��59�m7�6�s9�ԓ��U �D��y�u��Y�(�ܿ&�hL/��\}c�_�T�����(��r"�IȔ����.a��O����c�;/D 030Yr�r&��f���,Aۖ�IcV$ܙ����K��"�;$b��{S���:�)7Z�f?�+��l:��Z��T�d�����~�� QzKS���PG�8Z�2��# 8��>�,�ZD��gk-��ۚ4��Ս���P��G��)�����)����>��3�A� o2OS���G��Y���N��F2PDgT�[t!�h��q-����/���A�� �����,W�6vlF�7/s��v6� �R��
����϶/f���C/�'D���a]��y�����5��X�&VJS�� �����0n��I?�[{:Hw59�O���l[��ª▜�,�d-$�Oq�b��_��n&���f�B��M\?{� I˓'�SE�-sg��l�"::�#M������zhyP��"�����jh�^YJ���ɴKN	'�60)��h��l�W�)����?��ڱ�oDf�u���ysF�}��:�d��; A�b�:�t�|Ќ}r�M���#���&ۓ�6���j�hm��~���'�������;&1F�MA���Ƣ��o�e���C�jy'B!�ê=���$�����|t�V�T�{e�%�I�AN2��Z� ���������$����!��Bfyh��+��T��}ȉ�lѨF���dT�Nқ3��b�ҧR� �z^�� 8�`�j�S���ӱ��W�dIc!�w���cD�e����O \nA�O**�hö��w��$��i޹Zq�7
����<��^�3p+WH]��
;��q ���F̹�m������B`�*�a>��aU���$)$z����0��
�r������޴��8�R;��p""n�E��쾂�K�����"9߉��ʛ�Έ�PX-�.�G5��x������@�2*�5 )2ہ��]�S��gnߖlx�Wޔ;�)���U�����u�0 ]���2�%/�|vecB��M�m=}Xs��$\�xG�"�$��U���/O�mY�Y/�nS*P��<�'�Eg��}�N��)���9��Mk\��b3e�N��'P��0�b;��&���hR���J�N���Ы�����L��!�@Γ���Hr���i�+v<�DwÐ��oG���D_�b�@���@��V� L�׵��uT~��g��
��ZW	J�4���5j�<�|�WK��	;:�]�cmSo��+����c�o�=|�
[��{�Y���ZR��߯��赣�~a3H��o����)�}U�+fLŻ�Ĩ�6:������K�i�~[=�_�D����G�Jni�!�W=�{m��4�6$�?b��K\Jw���u�@1�`g� �M�Ie�=x�i;R���v�4^g���k�k���J
��ԅ~#4]樃�Ȯ~t���\�~��l�x-�Pe�k�&��Kd��r.X��-z2<�&����l$7�NGaK����ɜ�:k��7�����9����D�K���U�mr����x��ޯ�$�W~�*�[e�w����R�+�Y|(�t�Eut��fu3���ٸ�i^�S#3[�e�d~L��,�I�S�8�g�c6-y��J;i�2����l[q��c��{��f�S�ҟ�Ȓn�z���+����.A6U�ݱ	ܝHc+��.x�hb$�f��u]Mj���������"J�@{��I��Fn%~�|9=�.�'y ��a0"�@���B����ki<>��_<���0(�3�j'���8�;z�ܮ��tW���7��zВi�Ӝ��e��Hw�+ǵ}�lw�ܜ�>_O����^�#��jnY|�Ԩ�x=�LL*m�7
�>R!�=�|��! -d�r�X	nHY�<.H(!N��'����Ä���5M�ZTNQ.ih���]H9�C�|̓fT=�����2*V���"W�p�Y�� o^�ׅ�v^5Q�O3���t4^Ꮞ��
1��[��'��
O���vx]�k>�RB�P������G���8t�<F��������t�����{���������NJf� b31$�} $u��{S���(�ٴXaJ��ã���V#|ƁO��Ӝ"1���� ���[�;Ʒ-%��������o�95Ur�ΐhs.��UI�5XI`^�r	��25§�5�$nA���ZD�v��������GA{���MD"	�]�s��s�hM�Z�����N3�(-���>���)z��N2̗��4�-?�-��A��+B�%W��K�!��H)*0sa��k�����Աb�n�-���R�B ��-n&6�ñp)��.��A�S�y�qcƾ[c(w�@g}=��K���A�kJ�U>�" h2
Mx,����E�O����s�$d��j�Rns��At̫�j��-Ӿ!B�g6	��S�粊�X?k O���H�\�f%���qe��a��/�u ��[s��y�S�̳v�w�@���C�B��#O��o
��L�!�v����s�j�&�t���8O�m.^*���.�.N�g�����i�N{���&������;��KW�/N��x��g��5㱨/ˇpk�.�)���t�n]�V͕,\�Hye'- ڒ`o�^��}j8ww܍�1k�Y�g��� ˖�h5T��bs'� ��r����2��d�E��ԕ!�=�(��7!�	\-�$H�(�&�M�}���e�ц.�cx���͊V
;�=�k�^���EE/�����j���o_�=�'o˿�Ğ�(��@n,3'F�&9�̀���龉4ڥ�3�0\+��_� �����[��ù0iëEu\��uD}��R���kl� ��2���F����:]P23av��37*'���e���<Ia����(~9��@v?��IK���L,Ą�'l����丯�M��^E6�\�S'�P��e�֮�x�����惂��:�� �>����3yJ��^��[$�*i� �M���@��2
�f��J�{�vQN�o4��}[n ��q�\L�VD�26V$��k{��R/I)sd�j�?��}���
���1z�Iø'��;�y�]�͚������2v�R?84�1�e}�\ѭ��&'��Ϻ�ra�Hhk�iQ��+|<�1ݧ��n����N`i�Q�Kֹ��>�
��N�C���v��~�'W���<��9����?b��wH�U/�q*�tю��P[�'x�._��{�xҜ��߀]Ҋo��t����F�_��uE���^'�ѭ�<i��쳐�ʠ�莚�!�A�|�E�3?;��E���W�xK����	�'1f9-g��L�Y�䂪����Ў]߂�ٷ�f��;�Ӝ��>�����1=o�󭐎K�e,%�l�t�7��_��:�}wq���D��k*�B��\��������m�4� ;9/��y�Ӣ�R�<�V����Lʑ�9h�����{��`a�7wd��>�n�A[��������}��v�$1��3�i�í���g�lX��ڱ��"؂T�b�C�Բ6S#�	��f�k�.����V���*-�]��y��Zl`�I�	�3/�e�qW�1�c��&�R(�Θ��Ŏ|���B\��tw656���n�/\|x����cx��4?3�?E}&��]��CӢ�.L�P����P^t\�4@8�E�B9�bI�ɢ��K�'y���2^�3S�E��#dD���������ߟ�)�SB,Z�qҾEjǖI��v�a�3LE�iS��]"�I_it?s�2ӳ�������ݶ��0e̱I�����ëgN�۞�>'�&y�2}>f@#q1o>���}l���I�En�p���Sͷ�K d�d�_z��*�[j	U>^�����,~.��7��a���.>�پ�8�t�|�U�O�8�3C�2gX�$�ޏv�;�<���G!����(��ZX�� �ٙ��>��#�E��������Ѱy�N���Ig5T��?%����a,���l0+t��|�Wߍ8ײۺ��'���FI���9Y�/�����
�j}���;�(���$N���4֎��<��b-)a��}���ǱȦ*ԓ,�b7�D ��E�\S�7��F��=����V����pm��?V��r���ۥ@�W��G���!�q:��{͝d�T~�Ls&��4��(��ۻ u�P2��\���ON�
>^���é� vV+(n���y���D�͠��`�|"��U$o��XnT�^6ʡ��u[qЬ+��U����q���G�؀rriC��k�c2�� v{�`̳���؝�&��9B�t��G��pe�c�"�m��"L��=|���T\�)1�oj��#MXae4�~��H_��1.��ڤ���GA��'LVľ���1R\5h%�#Zg������6櫏����p�u�+S��Y@�0y���jd�N������'B��Ij౞��;W|�K&6Sd{$�ۺ����!ZΙp	%�`��z��*>0�`݌MA�,�.1�W`<T�L{F�+܏�.Ջ ����<Yx� ���N�O/�>�@ږ���RI��uk+Aܬ����)���m � :�ʰ�>nH�Wt@`��.~���_�ad��g+�7��q�VK�k�&ЌC�SZ�_ԺUtw�X-��T�5� ��K�U�y�ػ`�MgSi����.�i�٭�e}���-,l�à�܄N�t�h;ɞ�y�;��Ǻ϶�����\_9uwἒ>i�,l��&�����=���_���4F�&�R�XY�o�R^���1�� �6ʎ
����jfES��0���-��x?��%��������q���=o?R4t�������R�28��j����n���t��`Ȯe;�yp�jqI�*7 ��0x��뛎m*[dԍ=�n���O�<iO����j$�U����]�Kh p/�1��&2��d-r={訙1'� JQi����5�Q�ۙ����XlT�C���uAܴ�)��ԋ�$��oޅ5葽�q�0�ɧ��~E��虾�n�@#U܉W�{NZV�h�8���2�n]90�o!��%� 	�}��e_�v��s�	��:��3�Xq5��'�XŠ<�ׇ���n�v��X~?��Ѣw��go_���t�?���v�O;�9�?�pۘ��5H��wm�� ��L/
M����PR}��љ)^z��Kx0��M�F��+:�ȡ�*yK����Kl�(A��ҝ�����J�w��xjP�#����-FGl���X	@�����{������������+��O�n(�؝>������}�1���q����m�߰�gp%H5%u�O�h�l��wN�q�X��QD�B\���H7u�'YE��sx��J%�
L+,Xo�1bl��&��>����$eg��͑��y���`C��`�ȓp�S�Tqĭ=��/�z��Pw�3�T��1��%H����f{Ev�y?�̴�MtjLE"f���M���R�jTN퇗I.���~�{RG����D3���w�,%�8qq�,�u���W�
���@���4�YP�2�o��!3���y�0"���(��C. �y��'ުa�ʐ�F�ɂ.)���ii�:���	���ǈ���f�La��;���'��*���;�Ѳ���A�	5���l�<N`���z��zvة|l:�LK�M��*U��L����`��W���wx�K�uG�MCw���`���m�锠�d��`p�{�#�u��=�_�Ѫ!�1~��^��w�(ޛ�5�����n�U� S����c䠋�[i(�qNhׅ��FíT����������׹ؔ�C2������o��o��p��N�sԊ���)��:�"�_��ڲ^^�,��:\m}�˸�1�}��[Y�A��Z�:�'#`�$8M�ZG����(җi$�YdJ\wl����d��U�<���M�,�O������?5��Dz<�>�w�3cI��E0u�*��-�8LP�n
�imk;�b��i{�[��&,~�+>��
g�Jc��u��C�#�*H=��+���ʩ��
dJ�W'�</3��~\K���`Νz�Q�Ij&�?��y��')�WMKcZ0�U�]Yj	>7?�m�(�k��eO�AaRv�`��aV%3[�,z�:�� 
�'A<�
�� �ܐ�2��9� �����O�-�g0�2��<���n�滸��F?����}w� ���<ӡ!�J���Ö�8(I�?�+��	Y-�S��Ər�@hFe~�@������.���6d��%�GW3ry�����څ2�L��l�f���^�a�T��h[[[f.%=r{X$���X�`>���>�-Cgݟ�2p����vK�$��,��f��� ���n��%sBӃ��N�C�c��-���X��Z�^�Y�\p>�����)���d��`����sʄ�_�tBu�3�$ �M_2'9=������
���j�W��=_&�7�Z�"�f�������`���đM1(Dm�l3h�����+�*g3�3�*�!��u��Mq���Xf*�l`����b���SO3d�)�@ ��&\�54D��ˎ����'ȓ"@(��U�G�s5\)�f�H����O��8��e'���3V͟ݣU���<]|=,�e�'��}6�~��7�`�/,��Y���s6X�.l�=!~��j�*
G�p��,"��=�0R^\�;���v|�c�N�V��V�ɮf"�4M}$g>�LL"���P6
�3���6�"�|��ʬ'����<�<~�4sw����p�����ǨO(��`�� ��9h�K3
�_������t���'A�E�޵��.�aKZ��eo���OX�+�������_ǧE�_V٧JC���~d���$*�MT=��=��7��؃E^�D
�s�H�����'����-������D�����m�a`!	�5U#�������Wj���޽�jǒ���� w�����`J$������Xͣ��P�)��䩻^/%(�o����j,C�!v�d�G(=q�̜��í�}<�˱��!s⧤�sxxM,Q|K����*
����tm��MTmd��ڀ��1�_�4uG��uP% ou�?���Ly�j?H���H�P;�{k��C�6��B�S��O�l�6�B� 7L0����x������Tt&���ϻ���A�b����hp�r��r����̤;��܀I��בf���oU�����5z���G�,�����3D\�/K����Xλzi6�
��HP<�F;mq�V��b�����t{r+d���������`}u���7%բgU��p�j�Hw�f���0rK�����i6|��!�4zxu꘼���3q�Ǫ�I�ݚ����Jk8�FP��]/;槧�jr��~)~Bh�q��h��$�Q��+2(8���k�ם��^����*��P�C��.aT�ϙ��:
Ew��|�8����e�w��!bBk��T�������Y�5%��F���e �w��͌���1D>&:	�n1Sc�*��w�EL�������A���L�`;�&��5� ]�\��F�,�f�tk�3��Tn*�n���s,ݫ�L�U�Q5�Y�S+v���,7B�����0h=k�ŉ��]�MN��~˷���X��Ϛ�|�s�@q�jد�����H��ĭ�>,C�"iF�TW�d٧��a�K(��T�%�Ѓ�����p#RP7�JnWQʣ�_�x|0^w>�y��ɐb �
�#�D�P��|�yA;��N)���.a	�'iY*
� ���(5�)`T�#)��-�M�N�ϫ}�پ��n^d��.� �\����l�L�����G�H.�U�k�e@�LU��DMJE�}7w+����n�~thj�=n��۵�z�o|�?�|K.��7<VLV�a	�P8B�l?n�"���ʍ�
,ß��S�	_U�)�)��l�Ч�v��70R����HI��9�Ȥ�,��:��]�����sF�%۠6&`�b�0:W$5��C�FN�1}n(��]���|0#i�Q��ˡ&�xt�x�x��YhO��J��� V:�HƦ.}ohfu��o?��.b���>�.q�x�*�Dc5^dt&��2Mb�.`X�w���L��Q�(<�e�%`)�F�(��"jg���� $�$�TGLP��+DAިŸJϡ���s���iϩ�o�8Z}Np���%OX��
1~aվ��2j��C=<��ADx0C1{����|�xd~� �j��2���gW�F�PR$�w��QyC��)/���b�w��z���`㗦Cs;o@�̉�C�6��|�I�g�<~Z���ZJB�����5dL^ە��Q�9ar�b5�Kٵ<���?��<��z{%z�|�X��8	]���`g����~X���X�S!K���2��u���tD��Y�cx��Nh�f$B��L��c~�rtN��?;��ѐb˝hwj\��%8S����xyYF?6S(�f��v�!�X��>�D�d�Q0�ǐ�,�VK�*���|��)��dbUF��%�y+
in��fh=����s��u0R`<Z��鴮�w(����\��0�����XR���V�Ƞ�������l�Ů����OGQ�p-��<[�^A�R��׆H�����nK��3v��+�w;��c��G��2��oy�*�\���Ȯ��3*�_4=PG��_Ъ�E0������t���Z'�<gb�ZnU).x�f�M��MɅ��Ov�99�AD2�mW�J�<�kF(�Q��(��@;1�nk�r]c�Z��ۢ~ӗ��Q�J"����01�Z���TNV��!�NңGbܖ�[I�]�S�*/�>�3�p"��<�֖��|i���A�j� b��t}��-xuT!Y"�I���#��Pq��#cّ����6�x�n��mη#�+������X�>�yO�I� �o=���d�͘�s���t�X>x���w��af��������.U�����.������x�������,��؜�B?��^l��w"���Քъ�!׬�/��q-���[�a������ uf��t��ӗ�4��ԼD�5<T.����Ӂi[�L\^��B�C�K�c�a�|a�<��p&X��P"C$V%;�c#�gҷ�e�O�5&��rB_�=��=Tu��v/��pF»��R.��A�I¤$>$wE�vqLRa����εV&툍�(`�>|s�l�vt�ǅ?���c��;�_?������-�,��#�A���t�%�l��q~G`t8v��#:��ð��1�#!�}�;+6��I�2�zّd�?nv��� /��n�E��m����	`ٞ�NԐ�ʹ����%:0Y�?���JJ�_~��0z�xl�=gӜ�G�_��hs�����m/�q#^u�ff%�rx��@/ͺ���j4��(��N*�v�&"����mm_��*�ǐ�~��������0�Y�׏�5��͒�Z�_��Ɨ(<7�4j��m�
�_6�o��K39i v)��P���=�z��l"�c�z~�
G5���B���U4ϐ�o���U�Lr�t��~<&����gz������H�e8o�r��G��ڽCX�a/%�#w��(����
p�E���6��_� �2��uw�W)D(D|����Kk�������8�4b�����@�x��� �J�#���d�Z���)c8���Y]�	d�PY/ �
_R��L! JZ���WyF'�JФ:��>��E&�3]�F/��F���a�DJH��V-�3+A���M��{X~����LZ�,��k-�oE��'�7���D�լ�����e�/02�Q�n��ԁO���S�
���t�$����78v���,̲;ݿ;�ŷYj�pɻ�
�9���twʛ����#RYȸ|^5K�h��wh��ܬ;CT�7��\��N;ǜ��*�ی\;����Ε��s��a"�0+lҳY�Z��=/Mp)q�>FںtUn�����[|k�Z댲ҫ��ϰsA4����=�ܧi��^���J,�|�����w.i����!-�I �i��� ��:�W�(cT �Dj��Vc��7e(�&�
eI8���{~������
]������pѳ>B%�p�;LVi�"���t��$S�Bh���M��~ޜ�a��:z�7@��3�w'}���=�{:���H���j^�1`v-}�"j���Au�@@t� ����'��U_]�$z'ɦ�MWF�	���Ƨ�f�-l�_��̡H���f��i��*�t������S��nb�|�^d9�%vNp��H�a�E,��Kt�O����a|�TX�֩�e�V�O�&y!�<R��(�-g��/�\�.ZoW�,R,�����݃`lsd~���lh��W��T
�p��OU(D� ���])ԣ�ˊ��+���Box�p|^���^"Z7^F�D1�<fЊ:��so-������@�Aě����}�Je�rXp��mi�4zeD��v�m.�CO�:7 �!�g��-�|F,���<Z׺�#�G
Cש!�����j9,ŘI��zU�E�x���P�E𰂫"I%"3���@���M(ӂ�#���z"�6!�%�v�L���o����H��ge�Z*hL��B�h/ٺ��O�e����;e�i<f׽��u}.�J�8���\�0����j�����|̹4�Y�)6�]�-�m,䗯�"dXNc�ܞ��J�5iUͅ�zl��*��h�\�蕅� y]�ϭ�cZ�1:��1�>��'�!Uf?){�£�sB)L�҈��d�i��O�;vb�O4��&��w���%�TK�e�x������(�Mp��&Ӽ,P	[t��d����,�*�<*C��H'G��B������� �ә3��NQ�>�Ea��r��(o��2L�u��S����Cp��ٴo�T��o:�B��� �8LGe��{r�8��x�z�\�5��셳u�V�����(�j���k��~�2/0Om�6?Dhd�� Ę;���I��Ħ��]�u[$�*����*)�Oj֥U���a.WU_���0��O��7|�����k5�N���p�P]�Mo��s_T��蒞�.,���n�}ڏ���� ,��ʀ���ֱ��.7�iys
B� ��#����Ne�0S}G� j� �g���
��м�L;R��⚠-�'���p�3^�LIII��#�׸�'��z��*��s7�L���������55����'t$XE�e�1�^��l��"5G���[$��ѳG�G�f�/�˲s	�"���E}��)r��HGU}K:����h���K!��Udn������{���DFs�J}-D�7z���Iҷ�ah�@�����v+S|<���߁b�����l)�c�I�z������  �ǿ&X�]�l�Ke���E��5��U؍]8�he�R5�?�"~����0b��\}&x�FWGt���`)�������z����P�sX�^�Kۮv��X��DV��;�<D���-l�w�0f��x�GDu���_��ir��>�AZ��S��Z�{��w��t�Iw%`���@xB�.Z�T��H�c��9T�SM"��M����� d�ة����3�Ͻf� ��\m���#K�r�$+�����E�7��<���b�(�E��sr:�3߇{�
�v��b'��_4T�i����@E��BE6���%}��qG�^���BkeG~��k���q��j����j�zɒ���'�!\@>��˔�d�J�f�a$>���A)q�>C�FX���T�Д��oh����@� ̿�1y�ڋ1E�+=5���ل�Θ�~�'?~\�L� r�4�
�q%��_�c�y�c�^;���ҕ�L���s-s�ɶ�,VqQ8�V�(?���s�o��r�f�����**��>���� *E
q1D$�\��h��]R�-�+Bl��ހ�h$7��!@��ǹ��1�� ƿ����o볒�:Ϟ� ǩ�b����U���� 	z�6ƀ	V�N�%Pc�'�5桽���f!��M�A�=2����Q@�R�]���,R���~CE����b.{j�U%z<�o��04K���H�V�ȿluk`�R�ɝ��
����W�OAJ��
w�S�E 3mz���[�n$`h�ḂO��~�k�x*+�� /��Ktb檢����@�H�,�~�tť_� M3}��<s/�y�e�I�e���c 53�;�^q1��phЙ7錓�U�H!?��&�	��<\���E<,�^��������z�&[*���jh(�})9
K�_��P[v�u�~��g��\���o���a�{y%]��#��vY�����G�<6�_�x�?H��:t�Ϡ/
�6-�s?+3j�E�`yS��򪿙��kիb~�͒B�^�V�$Q#>\�9C&&���~b,|��bzb�M^�J�\����Ʒ�{,�j�[.(���~�X�Fs�El�- L����6&�r ����nK����g`��_�އ����z]WF���{U�!xQ��(K���)�N13�e�=��U�}t*e��ޫ��m�9n���DT"��5�NI(�V��4kJ�{� �����x���1���Mk.�3�i#
�M�������X;� ���y��fYI�5��yk���}`ot4�y`7��98�AD�����H� ���D'"M��2ZM�b���d�0�v�)$��6��@��L?W�қ�3�4���
�YΡ�FAwyf��+L��PON51R�]�k�����t~�{Ī��/w�y/"Sӱ������(٨�����S��c����z�W�\wRݛ�dq��
ƭd-��=����/zM�AiU2�Eid�=�� Be�C}Z.�d3(ҏf��5x���_.1�AMp�25�̮	)���$+OeD��蔵��3���j���]&��-���B��83����c*��F�w �MK����S�^��3���{e0��Y���\H����+1b���V(B����T:L5��Υ���-�d�Oj��$*ƥ�
���R��|v��0�? ø㾊��������yA��y�c<��M����3b�l� j��1��G���\@L�V���Ε3�h�r��({������g�׏�0]F�vN�Z	t�C�Vv�1�a�τ[�<|0y%}�ʗ��<X�B�����h����&�#��?5�K�H�ג��y}��� Hy5r�U�)���JJ�P$v¬ތ8/L��ò�̝V������x��!�e�����m8.\7U�r�7���z�g�����T�=
e{hm���J%��k���",?%;��EYS7���=@����-��!�n|��o�+�R�6R��|���#��7�5��Nzt��>/��S�� ���ADȾ;,Oơ�j}��u��f��K���oE��X�hy=���K�U�]V;s~	�B.p��E-���*]K��*�ıCu+ᰟ�H9]=	�t������<��V5��?��X�X��b�:�5N�Z	͙)Ū��e�i?%zS��K��k:�u�4r��7��#E1H������H*I���u�r�uK��¬�o}�|��@�9����BP/�z6<����,-��>=���N�x$p���n�.��uO�$��;|�����n�Tw@���i�G��ͬI2 �"8�6��8*M� �Y����]l��N3,}�y�#�ӷ�`�o�t����W�r��6�-�IV(I�� �tE6;R�c��q
H���<;�����k��@���(M�$R����v��T"�<5�Omb��!f��;wʩ�,y�'d��Y8*��rj��Kf��q|��c������c��J$�x�@w � ���'��fː��PP��δ�~���=��.b��S'I97o;���pgȇ�6�H�-ޗvI#A��5B��.��ɾ�@X9�1����"��:��K��-�+������C���8�¸eX[X��� �b��� � ~(W��0Yu�Y"n�W�ٸ�a�r��E�� ��@j#���n���ӄYi]��0قZh�@���dL��cp1�r�	ˑ��[�k���k(������C��՜8���o��`�����dGv���-Q@QgH��d�Н���ZH��shi4��t�n����/R�w��~�]9�q�+4��-gY�BT�:q�Isy2����Bm-�Ùy/�Vo�Jq�u�;:�=�4�*;$�J����a�r��7_�Y���S��1�'�+6�V�~=ܞ��[D�W��!��Sױ�S1����Eg-\�!ˎ;�q|��� ������mT����9��C���m��I��nL4q,�����C���g����)<��b"�9ԁ�Ӄ���+�Я=�MhG<���lIc�������y!���;���M�� ��C����tP�����4����N�-rm��Ն!�f��,?C(|�k�)�e�;�|���q�`��|�i0W+���t:7E��y��9�ɲp�W�C��ʻt�k�!��u 
���B��s��T�	VZ�5hS<0���Y~D�����+ɟ�3fr��MmV�\s�����Qo/�4�.%Z��7�n]���Z/f"֗c9�0.[I	)'�{�h�6�,˭�7@y*!M�B����7�u��/qW�6_����V~���F>�A��$�&�('�K���ȼ�_�f�쩎�w*�e)ƺwN�s���s��A�[�(S�2� ��j�y�)�
��pe�1&�[��/���z�u.�Ұ���ЮE0û��]a� ���Fa��V��
���ԉ2\�yShT�|}�Z_��Յ�礗"i�a��4���Xj<���e*W`��FZ�7Qy�yY��ƻu7�\��RZ����~.�$�៮J1s�'�p�N���	"��H�1D��8~k��v�(.������&�B#P�^aC��c�:'
�é�C���ѻ${�j�,�_�3<T�Anz�$��^�/������rku�-����Y�J��ۖF��*ε_��*���oߞ�������`�^��n�"|c�a��Y��O��~�l�G�靇�ɂL�g)���/W0</�;A��d(fG)FnK�g�W>N�8��O�Rӛ�;�.;1���vN~ke��K���0(�D�1S�����fzPRI�~���z<��������)�����gq��2������Q�4�3�X{�k"sf�k�^P@��w���>pAš��EVI�QÔ���1�u�D���j^\�`�0	?��{�u ����C����T���oS�!>�h�SnX�� �1>M��I/�=�U���;��#��B�	 �m�/ϵX��_X�9� ֻ���Hj��P��q���	�'���lk� ҵ�������E�$[B�أ��^�xw�� �9�垤V��ӫ�lI�V"�՞v�a	A�x��o	AN��Y+z�`���Wp�~'�y�WS�h����ꁧ�8�)H#�]^�SH��k���`�����y��<YKl;��s2*��u�Qn8��!�l$5 �TW	8X���Rr����Tٱ��[a����x�6	r,�S�/!$�:�W��Š�L��j����
 5���p�Scd|�$�\��BK�ؤ�M��ts�BY��֩T���õ�Eu�ϸ��(��i"^�v�i(��=�R������`�J�-��`P����y췺FbsS�l�V$�%�=58ݝj�ۿ�-�X�N��imIգ�o<4���x7$.�u�2G4u8��RB�}�sP��m�SiVR�χ����t�`�!�߾Ok ���5d�A��;R9C,UmG ��,�>\ U�%�d:��T������|I:{v,�+�M�]T\�Rh��y8DNG���l�O֓�=$u��?��YJ��LKU�π#� �Y q>*�A�x��)A�����b�L���
D)�[k���,�e	�A�*b5��,ޡ=���p� �7',������^<xA�v�m
�A�r��ܖ�b���Rg�!�� TA�{��-Eė��g�����Ħ�a"H�ϐS���q΁�&�u6�_9��B�˘Y��BVez=�qϫn�-�e!-k��Ss�>AHbz�d�!j�f�%�O���+�{ޤ�z�aD��[���H�B3��N����t9L[~;�kF��l�M{�|���|b� ���;<��}�����79����t�:�Z�� �ߴ�X�)j+�,��p�y�
�ս���,�>Y,+� d��s���f\�K���`�
�%��q����C��ѯ�@��:w���ɕ����8����d�~#��K���G�W)+�-�"��x�*(��@9+����q���(���c
s"�����Z .���DT�1�+���V��dߵ��~�9-�$)�p���k+9 5�����7�Bhdr;[�G���5g�#z���
x�4قm�6���+�ɉ�|s�>�~�
T\�]��`��O�S%	���6NGI���T{�n�����o�_��x�rɍQ:�S'S��+Q���t�@�$�_����d@�)��N����L��^���vM" k��9�g}�=5�'U��$�.ü���n.L(�μ)H�S�R}d���ʊ�E^�?��*�6��]�|i<�p��6�+6)m���|�xC��^|a�^����l����v�1I��Gd]�] �F�C�XkJ�Q�c����3>�c',�Ά���yj���S�4&�5��+��W�s1C�a:��S���.7�Y
� t�r���5ꌣ	S�����&*��yn&޺���,B<�	��BT̵%e���^j.��eq�-Tz��x��b�M����e�5_&�J�+�#]�?w(��S��� �w:��k���T�ie���QZ�9��VT�_z��g^�tw�# �.a�X#����h߇�u1��M�l�ZO��c�t�C�]ѢAÝ�=�IɩԖ�C������[p�ۦ�S�C�g�<�F��Q%�אC��L��r��9/<yqem6$�#�_#߽w�C��o��D�H3��2�_<6���
w2�qT�.�u�A�Y���ʩN�B�]t$rV�W�sB��Z�-��M�K.OF�I��H��Yu�"w�rȻ�d��
�?�ϵ.�#X��kp�]4�9-�V#���C��~�=Z �vW����8([�8�.c��\9��V�o����O%t�ǋڦHB�ɀ�2b�KV��)>�Z$9�o���z ב0�_
��R U�f{�.w���~@/�C�$�K�'H�(�G���@O��tS�L��fo>�P�:� �N/��r6��Y�^l��ۍ� `,�־9��\��{V�����+��;�YqO�BZКl�II��E���[�{]P�����:Al������\��u�_��[��{C|;3������P���O�>�:&�����j��mys���2l��񸺼.��*)�&���ۈ3�!�_�6�B�^ӡLI�[���^�K��#��T����_��};���h�@���P�^�l��\��X�9?��i�fS�5.o^6�A��|w]M/�iWG�:%/�LND��U�)������۝���+︟F����|�f��B����0i��'��\��tF�h��XԖ�V�/yϋV亃5���4�R���_ӛ���b�!]�P�q����� ƿϫ"ű��Iͫ$PӑE�+T���p��GHI��w���gV	]�	&g�����]v��U)~��)���z���vh�L-nw/ 
A{��z��î���w�����Wf�����b�c����������p�=Ԫ�4J�U]��%�	�����!�o3��Ѕ�2d�C�����ɲf��y�N��M�L���_��k*EX{�|^
t�Ʀ��(�"6�RH�����C��(VtQ�{A�q��A�Hy�6���Y]�2�x���g�/��Ñ%���z�� E�ɈЩ�@Y+Ȣ4�y�b�L���_*�aC�IC�%�£�_�F�=ݨ��ꮈ�0�`u���e�Qts���K��3x -�n���)J5�<�K�w�]��X�n~[q��L��m�`�e�F�^���*�|hA��w��K/$GƮG-��0@�>R��Sn�Z�@p�<2���{#�RO���ܹ���Ig>����oHk��o���w�;.�e	�]Hs^��n�p���)�] ��c� k _��@�~�J}����<�-Hj�x�I�@�(%�/���rV�{���ȷ����
�GS+�`�T	��;�E��N�P��Hg�A+�Y��,l�fS �4��H'��Hg������K�hn>�Nɛ|z3���f�Sz�ësͯ�a���,@�_��y��ªN��C�W��e�D��@� W��,��G* ��~Om13���1�Su3��vi*�󤇃��8����Z�QZ�>��1�e�?;�i�١2����<�U!�,yS�8���DOch\��8g8��Q�93�?��#�u8�,[�ol/��("�ot��w�z�4#���R�ǎ��A���cJ�p�:�g�u�u���fs���>�~��^7v�87Cۅ�VQ�ǆA�����T��'0�ZG�S�E�#lw�"x�����V�(�OD�͎m���Y���C�g/eU����'����u����pޠ�^S�1*��ۂ{��ĭo��ٜjc�E��>E��U26rQ�+]��?�zh�M�0���85P������e��4TĚ��5{)�\/���ƨ�Cf��߁������
x��4J�ʸ���Hv+݌l�/���Ɠp �J<U;5, ��XG�ab��`��Br\y����zt���i��Ey�E00�Z�c��a��߼A��5j%�;x����p6���@Tߌ/ɳ������RkSm��$|��6gta.��ǯ^ح���ڣ�4Z��3( ��Q�u�}��'���
�̌I3[k[�=ɟ'��^{�5*�q�J�]�[��Mo�Z���w�������2�N%��_�kS�4�{3x�(�:a�/B�+|�ۓc&�ˤ"�G���������&Zg�e�|&GvsL'�y��4��4�\A�4Vʺ1Rk�E2�N�N�}��RvU���%�D�N<1�f _Eg�F��@�^���Rݕ�G8$�۵��۟6�RvJ���:{����O�/�q"8�K����b��b|Y��ٞ�qy�4�G2�+>h��q�v0|7J5H������҈�0i|�Q^�w	�ZԌ �(��Dxzw��q����M�>�J��Ю.ӂڇ�tkj�lZ�ul�����t9��􈻍�I��!л���8�쯛��Q��p��a�����O��Y��Pj[�=�:�,6;���}��O�_L�K
�%�|G�mc� \�f�[��r�+�����PZ�e�};K���B����pAIc�;y�H��Y��ppb�*#��t༣�6mX)��SJ%�h�d�#����;�֭�m��9¥����@g����o}0dj��R4����F��#80�V �:�������}l��CQ���ȸzٻ�������LבU�3ա����Q8v�T�p�#Q\�s��� ^f� ������U(�/��Y�-l??�!fjپ�ܰ�#|c����Y4��Ւ_L�	#v��`�-2L�8���nw5�.��*�����n�;����;m��w�V�yn�:�gY�x���KuAѼ֌xܰ;��Vwe�v�5Y�E��1����&i����|+�~/ٖ.����ChZߠ)(��<�ַ���X�	(�/�n`ܭ�~W�0��A���,=M�+{��^t50��1�M#_0��"�<ܩ�z���3̺x<R�:6�z
����~�ݟ�*�*��@p�#�f�*�նb7���Yq-��~\�N"�ǟM<�2���m;����
t;cJ��S�^ M�.wB�θ���)��T�E���N����O1Zr�j_��XM�QO�⪳���c�{�i�a���rE�K��q�A�+��r�;z���~��P;W�i?Ɠ���3ĝKxM�ncG�ƹ(�0�Ai������
g�7yQ,�`�M����sP�s�y�M �,��9��g� �jSa��U�mr���	�;��~=Ғ7f븡W��!XG!����NJ�iv�V���enФ�n!�1�eю���!��Zj/oA7���kB@�?����Ӏ3�6��~�>��]ﻏ !#(�Xz~���
�.1�����1�4�ȍ�^+��!7@��L��7b]�}i`dU.��m�V��(`������>YKD<}���R5T��z��oK��.����Zp�0]�&#t-Nε�RS5�:lQ碑�s�,�=��O>�mE�}i��Bc)�[����VE{VTNKq�]�p`��m���;�l/�:ӧKɐ^{��V�~r'H��֧���W*�7wT���n�m���.�����M���v���_C?3iA�MT9�%]�@I��azT��+U���M�����b]j.��j���ԓ8M���e��U݁�4��_G���\k{˨�6h6d�>+�+��a����e:��&ɥߜ
��,��Q&�UV��Q�q��a�����$�S����.ՠ��m��6WF�\�*v9��s��>���.`} a��e����95���Ӥ;d��y*��,�:�JAf7��O(_�G�Ge���آbĴ�jL`1�G�R"\B(j�?�u�/Ih��쎢�gܵ�U5�._�{&p����c��Aj�~{��VwbO�S�����ӭ��n[���{di ��A��F��wjgCKB���H`��+��%vof;�a��[��ڲ�vhP����C����\��+�3��sq��������'�g���	@�i,@^�Xl�O�s�Rhȯ���1^�
?C.��Ǣ���Ȇ��7��W`.��S�7��L�K�������������K�MPly�7���VA~����]lǱ&vw_9�� ��=�����x�H��d�[+��?=�{�|S�����M|Sq=k	�9�?�{�B&-I���9��9��-q����T�P�B�ٹM=� ��n\���g8�6&+�~�g�{���j��?ί �����p{¾�>�$�5h{�H��aZ¹�V���k�l�|��6�Z��(U�뇠m�'b9����$ǋ�:�t�lH��rI��2����%�8�+`$30�x�����2L<8�����4���8�p���sӟF&�*�����Ì�g�'�\�IV�	���C�_@#�nH��iŨ�~��>��V�9��� ���z���Ҍ�y;�f�f� uB�Ɠ�M1yE���NĿTwl�4�zSSV��	N��ʛ����^CU�ǣ5+��d�E@��8-��5SDJ�$/�{^۹��{-�eO��j[U����{r�	}���&�n�#�
x��œ�P��{{�V��oUcr�S�*���F‼���?76���Ec�st{�61m����ܖ�a��:<��SQ�$�	�������U�����-��E��F�� 2?�,K��ue��Ր�e�ם}{(H�*���ѤA1#���od#3(�Q���?7��&��O�Y�'�7�JCE�ap�􅺮��}�N`�?�D<k\����Bm6g��@��� e4k��݀�a�vrz�u��ɘ;v��5`��U3Z��5�I�6L��bO��\����0F��x�u(��N�9�%�X�$!jxTo���i��nuV�]M�f�,��<]����3�f�`w�E�)��W�dKKp"���U���]�z��R&�:�`���Ч[r{�/��*JZ9� Ff��x��s�j��K�/0��+��˼T]K�*
��@����)�&H�X�m����jZk�/�ɐ8Ph(�F]���]�ָ�Kȫ�{����#��}���n&E��b%�qY��R[���li�@UԆk��R�q/
,"��귕�ϫS�� e)>��@�]n�����USa2v���u��)¸�5�5?�#���Y\�a((��j ��a�fE'<��c�����%����;��e&C��K�l��g'Ul��u����"2��f8Ym�oԚ�:�eq��(�{UFX����0Z�dw�՛�Q��z&"�*������p(	�¼, �-}gJ��C�׼�"ߌBq!����ք)������&�t�p���A�PVUE�H�X-��7n	2׭1l��/�!�/є��5�qQ-��)����bЍ���f�EY��6:Z��r��� ZX@���A�M��ь2>�1Nu|�*Kg���4�O6�"�gZ��4D~2���%Q��:���P�`|�[�_����"��(cW����2&�g���H{39ʌ$MQD��y�~y���Ɲl�1ؚ+��!Q�ݍ��=.dx8Fw�2B �=�Р(��^D9��r�n���0{c��f�t��<UU�eӕ����8&�B��rL��F�`�V�՝�*��/)�eV� ��A���g��i����P��OJ��"Ҡ6�!�29�صi�E��&�Լ���� �KRl��3��x�w��&la�GO�>���:z�(�}��cG��`;��k�����a�${�q䁅��c�[j~��1XT{d����s1�m�W�\ES�7C!Ʈ��S�pa��