��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)��<�=�!ʢ+���#x��ȴ�jo\vc�l����0�*E҈�u|d5���EW(SصL7�/��A���1n�;M��%ڊ�C*�q�$g��=����S\$+R=f>�ec�^�=;d5�:V����)4���R����Q��ߠ2?�L��ɯ�B�Hߗ��[�3x�����<��y���Gz����E�5[ �4�j2]��&~6�iK����7g�5ʓu�a9�Ңp��.$��Azgq˸��.E�b�w�3�`��CF��U�̓V,<��3���m��M��u���c���J��bo��e%��т�4�A3F��wc�g��F��M��6\�`�8P���eT7�4������~�Z|��Zd02���\�M,!��pt
N�q =�;��wK������~��O_)~|�d#��x�����9;[�Bf�6��-r�C�*-�j}q��Tmz���������z?.������J��xE.#D�"��;��yO>�w�K@������-#�e����z�n�*x�*0�������9��R�<����ۥqd9}@�}d�(��O�os�����[�"��)��G�I7���;KgB���^~�k�q?�|�x^+���bb�֟��C�>���S�,�|�dvu7D��՜���:hs@
<t�������8�EeV����X��j�B�p1���EWr���	G��������W!�3
X�Z?��s�G�K�_-�& c̔��X���ܵ�MfW��Eq�p����֔�;�tk 2�O����82I͚��=`��k�K���R��6X�q�\��]@k����Z�21ց���2i���[]<� q)��'Yo!�s���#K
��I{
��P�UÖ�[)�I���|�Jυ�6��`X��9�Ⲕ�9��æ�H�g��ά���>U�0�|5�g�r)�ɓ=�Hظ��H:!4N^4��f
�}�2Q�KeW���ty?��[|��T�.�Tj2�
oI�s��ȧ���"Tw��O����	��q
[���T�E�����X\�Km֎�mK}W�32ZT��0$���]�PS/�M�b?qQ)�=Qrmݭ_.�'m�Z�|��Ak��zdl��m�D$`@'`�M�H�c7�Gyk�d�Nzݣ߅�w0�Ԫ���R��_�8����QdR�A�U虺o%����!�����j�ob���K��Rɍ'�)$h>A���y1�a�.9�����;7��-�hM'��^è��9��A`ۂ=<(�37	V[+�U�jx�!z_�*l�O�o2�k�l��������8
KT|���N ���������r������~N{�Ji7ji#w2DM�,p������<���G@�vB*f�\!�2o`��I��.1��gV\�M�&0��x3e<>��ܦ`�N��E��w�G�7ckPfF
C�E%w�ڄ�+8E��?�/�uI�@�1me��^^W�f�(��5��1�\�a/۞�y�I%L]�
\�[֣�&�d���v��z���9�?'�_K��W��-f���L�F��N��[]�*p��@�t��wv_�f|Tq�p6�݃m���rL�,B�M�s/��n�1:���^=v�ĥ���!s��~��Zو+J}��6�,�ܿl=�&����YQ$il26 O���I4�^jj�9�R
dl
�=�uDc�m�G����ɪđ�Z_q�3�4�T8�q��T犕�>��+|�@l�J�����ھޒwi-�� ��mśB�g�θ���^�&Lx���2ě	t�qm�J�*�Ҭ��D���*2�,�δ��Hvv���D�)\B�RJ���WS�F�ԇ%A��L��%��j�6�z��|��D�e$��rYJBWfV�J� ��θ���A�i^�
���!���e��I�~��:i�Č��=�X��^)��'�+�..8�d�`Ǯ1�yu`�n��_�_/�(@S�P:��d��p��O�#U���aC�c��N�j��+MB��x�Qlkվ�>���R�.X</�a-z�%�m2��x�*�7}YR:d���/d?��č>��.�
E	�[���N���y��?���"��9:�J(��� 	�MuV�2��}���Q�禛���N�D7<�v'�B�d%�㣑`SA��Ψ���+�=N��W��Y�4�ιh@��O�C'&�{��F�G��5�����'�t(�}֯���/�*�w.�YU�D�}h��-��)��� �Ʉ,-mf����<��)�h�W�O���0���|��;�_�WUNjE�0�����3���A�6�\i�GY�r���&I)���[u��܎�]�s�vxa�yY�t/FC%{_�!`j�B6�27x�kN.���Ee�fąj#��vP�?���w�;1�ߏp��Y�Q֦�G��N��n�6�g�,��H�D:���2��]Pg�S�fd����TF�x��m��@�Goc�+�,�p[��� U�"Ţ�VM�R=_;v��3�󾏲�^у	`���|�T<�R�:�s��d<�/�`Z�q]Qg�b�2_�v_e�4|K���	F/�3����f�6ŝ��@�5]�x�����8H�}w��k���M�\i��vEZ/���q+���/]���Պ>D��޼H���Z~�5M#l��`a�I�����2�*ZP}�xh�I3�2,��n��i���������J�
Uan�;��˛�:�+��<���z�P�ȅ~��[�^1g0߼8/����h�~��P�%��]��
�0��x������;n������p&(���O���@���9dCF��֩�?+���yq����]��W��:j���>Y5~>	:��л�F�q�%r'�8oj�㚬e]��:�G��v��c'4i.z�����*aǦ�e=��]d �
	\X�*�(hpɒD>S�����d\��EL���:�o�o�x�-��E]������_�+"� �5����Y��� #r��pϠ?�:8#�������G�5YC�rΤ���dk�7����8���9ٌ#H�e���5�3�u�ŴڎU|W�/��OP�B`��6�k/�T�Fk���++2�lK�*�a�5��m(ֵ�&J���H(#��p�aM�ՔK�ȇ)�Z�wÄ6/0CP�Z>�4���3/�-8�`*AF�2/�*@�C�>kF"���Ԕ��E<=%�9��ϧb
ٺ�r5�� e�;:��8��c��ܑͣ���k��p��A��vP��Đ;�eV��-�3�	E�l+2����;Ȩ>�!���_@ˡ��f"]t[Pڸv �J[�;¾��^��}��N'��VO��&������b�� x8�:$�郇%����IɌ�T�&�G<Y���@�%6#��� jӽI:\�L���cgxv��e�Xto"��h��1?��:����KS�&�c�62M<����_8�Ӿ�f?U�Z�H�j�eQ���AS!*'B��6!�����N��]#*���-���A2��L40�کx�Z��21�dc���*$h��Sه!:%�"��Rtހn�<M�Sz�D]�}�z�*�������7��T�q��χ���E�V�x��VȪ�}�_�B)9�jF��[n�
�V&��5���XZ��,�g|. �<�i�KK�F������t�]��xW�c-���j�V��]n���w
���I�jO��F���6�,�UK�ex��ug;��}���*�	��#N�@����H��P}�3G��%�e��˲�X��*@�L.�a�Oe���� �s���RL�f�Bp��$�,�N��;\�r���u�:<��)\���2�j�-��~a�$p*=E���ǹ����S���N�0M%�ji�glW���t��2�D�s7<iRo�-�u{ʇ�
�H
�_��
��z[u�pD���b���ċ�J�̈́�*��ab�02pw�Di.S�t��g�B�f���\����0���^�]��hť*��;�!�<Q�a�!K�%��weB�R��XnL��*y$J�V���Xr��M/d���j	��J�*[�a%]��/|�v���©ӧ쓼��R�ȋrħ&�����-@��T=\'H�!��F_5x�|8r�|��ë�,�:*��N.D�ވ#I�7���ak�1�O�V:7���W�z�|F����V{�pH�O�=}[9t��/�0��E��%;����l��pY�*��vM�;���9�_`{��}ʚ�t�ංi�H�1����|�	ߩGȮL}�������\%iE��VW���Gk�2�an���*G�����9��UO�^�,�W�nS�s����
���B(�.�\ C.>��ls�,�km�����+Ѹ���Y�(&��~y6H&�����I1�z�,�r�����FZ�S+ۿP�RB`�̈]&�{��ݗ��kp�A��W��Cr�^[_��W��k�͇��e[��G2��T�L�Q���'��W�i�evu�A��W��K D��-�=EJ>.��.D� Hw:�&��_z������l@�2�g�^���u[�*qs��c��K���3Vg��a�$���C>��4�ҭ�l��;�� 	�#&d����%Z��OK�&ț(b���f�^�������R��?���>��F#�%I�K�a�y�n�fP�ZP@lu��_Q��O0�7�l��[~V�Yo��Nޘ����$ɨ�)c_,%4�� �헎�Lt�h%p���V��XUK���e=��h�5���I.�Fyr��l�ڸ�[����l��a ��ї1
\�KBq��E3��gi9���m9'�*�4"�T��	n�K�p]�R?T��O�S�'���:��(7"�j}�Z��;kS��O͡����YQ��.���Խ���'T�-�y�`h��OE:{�tI�+F���H�?���Ū =�^�%���rQL�+G�w	U�9|�곧3��_�G·7�����9 1>�m�P��#��yٸ�X��M,l'�����%o6��M���K�\�����F���G ��`�bj��	���渡�{�T�"�� ؐ�R����_��O��Q��M��X�Bj���wb���v��kL��lT�4ދЃ��4G�h�L��e�ƥ5s�3�t�Z�P����"_��4�v3"K�Ii,[�t(G�#�,�����xh(�ȿ��_��'���&���N��!�z�KNЦL��ѣ'�j�)�E�y3���`_�ٯ\a�۽�b�����=���$�ڹo-4  ���IsR�p�f�_��nF �(~��|6�Eh�	�{a咞�n�W,A-@;�^�X�" ���#�(��B}��k=k��6������� ���	7#�!^Ύ�zFi6����/>��8p�c���L ���O���ŌT����),1����%���X�F!E�:8�P��1o6��D�V\�ы�w?c�=�b5%/�4���(�|�O[�.c�O\8�!��Ry��LY"@�*�;�j��ǡ���~}6�G��_�{3}d�m�3�n���E]]ރ�;�jS����+��w�̴B��{�VXD���6w(<*,�.ڧf�wg���/��q�b������I��L@29��a7�5�ÂKƺ^��X��kW;�V�M��E��hDp"�=�~c�������`o�=NǢc��1/��o3 `��r��b�6��M��NB���I��c��U@O@�5%R�C�x6t4*��ӇS����= �� �% w\m{����u$,H���S�HA�ǀ���FC�SE��~,�J.���\��1*^��m�EuO�x�JqmҸ���R0=~��f�%5H�VDfݚ�>���m�*[��ɲ&wߎd«N�����a`&�(k�ֶ�^�SM�8OOj��ɷ.���ǝ#�2h�����u�3[SwnզGs"�o�.@�DT
V�h��r�ȏUA��T�/B��u,ȋ��W���GZsL���1�/�T�;��S�ͷ�:�@&1�WZ:΃��@�a�b!4�֠�e�;�ej���U�^3��=�Cd2z�X�5���sCFl�ؠ��Nݑ�ēx37Haƨ2U�2)q	��tUY�|?@Mop(MH�<���%��EY���)T`��8\�'�*�2O7q�ˉ�"����!�
���
#�$�dF�l�N�b���$�k����tpS��g{�3��'F��׊�;^�W�pS�a��ބb��EQ���d�w(��Ƙ041��Ay���$��w�����O�l��(�h�'�	���wY�o��\$5c$���9>hϼ��O�*����>���r=�0�Q;����@��8�;�9!��:����34��8�0m@�2f��IO���9���x�#�>(�U �'��&b�4E+O2�����<Dt���'cl��"!�5��+s��g1��Nk��u��+���ĵ��?#����s(�0� 	��<V�Gc헟L��.�'�����}L��Ii�;7�1��ck�7�d_Dluv+��W|ˁ�[4��8[ŎZ �_�{����uҘl�f�!M�k��_��WW�G#|�5��g���H]Fnaɕԯ&��cD��,]f@����D�,;�|дS���Ŋ��-Շ�L�-$�V�N�r�*k�Ԩ. ���h>���<7��d�L����(v��C���K-�6�*��0�s�7�	�Z�Mj�,'���W惯�O|��{SC��mcu`3C�z��)�u�Ў!r2Y��Eu�S*��<;o{�~h����s�s�=-��&��Q����p�T�-��aK�-�ߔ �H{t�!n�J�>.���X ]Ħ�u͘ޮ�kPJ���P�9�F:@D��r3N����1��7�Ѓ"�;��!�����Tla��mf�|P��n�Pv�4]��G%�����M�43�Ӄ�6e0�e�V,Q8�,i�6�Q߫����>P���]�񿧞d鐻hC�Ua"�w=��i�f�IB\1:�f��v����w��S[V/�
�m�tv�d���8*��-Y�w�ݕ�Q����(�_��-]�=���'T�{%O��>"����p��lFi��������\�%L0�D��&�~B5|Z
��B�:�P��F:�#vm:Z
�@�_�.|U5��3�fF���,ejoy��V�f�6���	p�]�;�S��SKC�,�wh?G�m���*r�F�q=�ޓ;+�NH�q��to6�z�ً�t$�� ���f���a{ �4l!�}KZ
4`e ���<2�f�ξ��iy���lk_sa"�1��昵�_K#Cy"�ˁ�\��w��k2ʵ4��H杛[}P/�R��z�q�p��J�dl�mݵg#�G�`Ȋ.ز�]b�Ou���e�>�Q�R� �6&a��8�;�� $X4���xa�S]/m���<��sH>_��H6��<4J���-Ot�A�k�k#�(?�"�.FKw��-ᴟ��NLڗD�nl._�= !y���U����y俪f`���\������y�ۻ`����yDkAa�s7`͞�*���d�)���_.𗨡���N��R��q��H'���g�:t�B8@-]�$Qv���^� ިE�v�?ܖa�7Z�R�]�{���,2�J�b��������¿��\$@#�;�3K4Ȁ�Z�)���ci&,x�.�cR����MǂKh@�x8��<��~I�T���X� ~-�J&��TfP�B��i? �=��%�>�C����c4}���i=	6��>�|�)ھWQ�9k���aH�P�l�s��r��aء�c;��4�O=�� &ˍ(@��+W�7�7��1�ʉ��׋7��?@x���A�ܚ�nQ��u�����"��JL�A��-Չ�}7<4s<#�?,.�ja!�!��8���+��m.�+��1�� Ug+�tٰOڴb$՜��)��;xD�R����7�#���ŉ�
�7S���zy=�3�.7���Ӆḅf�(Z+����m����#�#���-LRD����*/L@�=���;���~��w�4-�x�Kg�_��WYPے5e9zat�����ǋy�M*~�W��O�#�v�e��[�G|�f��l�vتUOI�p7��8Z����+�'������5����z��D[��f��,~���V�9�~(�@����*��ra���Ý��8vR�Hl�Cr�t�E�߶{��Tތ,�Nt혅n�JW%�'ԗC+�S2R[K��P^1�|zjvl�@���22v�E�s�J�F��BV�:
D��=.���]�DHC��8/#ztC��j��܇F�d��y,�.ԙK��0�?C�R�*t�pǖ�dV=	�s�y�w������ˢ(�F�(G�z�CƊ�vY� \�f�n2j���G2ؖ�������}�
�M�
��vv���] ?|œ`J<��G�]�*�}?�	ԀH2�h����	�nFd��{��;+���C4U�u�������4g�qdo��qG*V��	+��>�,MC�e������H��*�����R�b��p�������;����i,��j��.l�A�֪������a���S�ڡ�K*\��}R3�5�����?���H���bQ�N_Wf2��m8�jH��˾��$��x2o�,�n�z�w5	�`�����b3���"&m/���9t���S��-�&3P3a�b�n!��`������e�����/�yW$���TYs9�ܰ&��q~1�)��<��]w�xh�?��1��Z��P�.mk-:�[���Q���v���c��A��+x0�jO�|��"� +�J��-�CZ@`���q~O_�Z���{B<�ű"���H�Fr<���^+��(�S�p�)���}2=�B�p�*���Rj����e��(֜�����|+>�[���w�v��Ώ��{[ٍܹ����V�Ss���G�.>Ә4/�\`�#GED3	����nBo�OOa/��c�jJ]����k?��D����ӱ!����1T�@V��=�M�ˍ��+��۹�ߚKڊ`G��Kr{�M⪭tz"*�q�\�Ɉe)̲�������/O:�@t��������ǰ�q� b��R��]U���J�6k�BTԡ1SP
&p��*Z(,�^6��P���z||���?�7��5��a�@G��*&�3p��]I\��&�n��gt��ª��m��ڵ�A�w���T�)��� ������k���p�F$�<4��"��K�YPW��|��������x�x���9�9�s�/p�x�A��t�G|y�I�Z��O����A�jO�6%E�q�}=����wq��V���QH{i�!��|5�����Q-��sl�|�����Y��l��6���6�HS�$̂��J�=��#r-x�,[c��!�j.	Q�с�G1����Cs�+D1d�#:c��x�����l��h���+?�@���==��W��4����z�d����.�(Up�����X�|
1fl�s��Z�ks��� ��A�ﬃ�r��#<� ǽ�.X�"���j�(�98���ϑI�Y��m�
Q"%Ҋ�?��Yh��j �>,��i���x3SW�:񊱅hԷ$h��ےbJr�G��m����z�G8�����j����*���_\rͣ�qu�8��������|�ƶ��ϒm}�o�*#�d���۸���e+�Ǽ,,���E�@�b{�x}�k$k� d��}����FI����,Z�tS�\���D�˫��������<	.���xp(׉��4�tO�J�g��C��aLd4�,�e�9a���(�fc뾴sS��WP�X�a�-�T����jܨ*;�û��YM��������g ���Ǆ&�����"=�9p<gvm�n�Foci7r�},��|EE��d���y���C:�}��T�������]��OGg2ƠA�D-�ت���?')N^����Z{%>���_u
}���G��a������6lQ6bsq(z���$�F�.V�
I�2�cT���)��C��-ތ ��|����QH��hj������6�]M��[6$F�~��d���f&`��#���/)�<�^C{�_�D�~��Vf��i���@�sXG�HB�'<����k��U[O0 
ΐ�H�����A\�=��}��	7zg�|�6m��lJ1�ѐ�'L(�򐬜MS�	�"��.I�
U_�D�K`�c�u��+|�L�.��:��M6��N���ïtkЛ�d!�����AiL��P`?ב5� vj�7b�"ܯ`�/�&E���kF4،�7�,m��L�n9(e��@]/��)n���*���_ϰ�gfo� �G
5H<�d;*~�jA�c�)�>�3�]�+y�?�/I1H�V�����(s%��$d��y���|n{\�mM�P�9h����48��>�96"�M[&�43�p��L9����x�gE�{��ℚvn#v���A�1�b�EG;6LN��X։���ǘ\L�u�J�,���(mHJ��m���^ ���+�AL���x��K2��X���&���`5����X�(�uK#ݟ���ړ�Ѯ/�<nmN�����3E��3w�.5���NڜR�
�5UO�1�G��%�?xu��M�Ҵ�X~0�+)�nny��{���f�|�j�5;�%T�!���{���·���
N����R<���>M��Byݗ�n�z����`��%T�æ��P
x]8����nn�	մM|{�X���U�U�����韜d��I�'�a9QF��w�3lB�H�t~��r��A�������6��93_5�p�)+��!4�ǽ�"���E����^��ӗ�����ǁ�u*͋\��׳��jJ�bI!ᙀih#S���8[�~��q�@��lz2�[(�N��ҋ5uz�|H��Z��g0��.�*���ZS��B��=^ _�S�z��C�p�X����E�$/{����4�Drʁ��,��31J�E�p`oC7f��oR}O.�x~���%+a�cr߈1�����ƜH��tn�Y��ETX5�ڤo4����Ah?�'i`vR�П�m��'��4�US4�*F(�\w�� u��kk�����5iBqT�T]ڧ�w���h�FLC�/��~a%�ߒX%�N��c�ڙ&��a��M�$Df!
�B~WJ��λ;_Dw��ߔ�����|lg�զsI���M�/r�C���������9�XJ��?��Зhd@�_[���bx��#.)Q2O�8a��H�hնk�p�0�lO������+eV*f��o�S�hd׻�D	�7ȹ��4�K�!�*���V�ˣ�d����ϗ�L����4\�Ժ���s]<�*+��o���.@�B�o����F"�k.�- j��t�53`YR�� �K���bɍ�� ��]�}�3b��6X�W6`�B�sl�u���xaQ^a���
u�B���wLp3��2��)1���O�M�C��*���bʨ�� ^�S���Bi�9��7ӕ`:�#����BԘnS��i�����	�4�,�wOJ�Zy۩���R]R�����䕤(M:�Q���߬��8b�����]�e@o�Y���>妽�Hx��vMݽ��?�N���]�;�D��2�Xur��v�yd���	���������4eQ�#G2��H}6�/��H���Z����\bn��聠Sσ��ìH��T��,B�d9�[�.��9v��s��?�� @n�LE���
�0�������F;R�q��Dƙ�$WؓEr�?q��Tq�����5X�B����`I3scV�j3\�ۆ,Q	['+�	�G��p"�=Y:N���E0U�	Nh4�h*�8}Y���#�]�{�6�2�h��*�	GA~� &�ha�4+�9ŭ�du�Bs�p_���YͺC�#PM�~�%2��隭�c�����"��X�M���`M�vD��{4��������ϙ����o�\�1�˄ ���͗�o9}9��!����z�ˮ	�y�����y�lHb�ml���.	؅��*��mc�Ʊq�nC� ��E.5Q}a�˜�T黀���ЏI���hU�3��D��u�P�V��`s8X��M[�i�M;/�eř3��2UJF��X�gu	�vo�AߜU�i��Z�g?h��q"�ʾ ix���S\��:�O�)w����[b�Vy��x���\�	y�������dw���� �)h�-fw���$�^J�3ML+�}62�	�(�7�V=����.�{/�z��޷2���AfYi�U�S��H��99��
��_Gqyb�6Z=�v����u�[.�\��cM.�}�
t���ק��%��>mW��%��]��L����G�]5�<G�틫Ve�#5pk��g8����Zp
vu-<�q
-%g�P߮�]uM��@/=d�q� ��:�H.��E�()�e�)����,;a4iʂّ�r�ó<&�\��C#��y��a���o�R�
P�AK&��M36,�ŝ�\�j4��80���`̥�}�}����R�w���^����C������M����|9��t�鬪ȋL�S�\3x�K���`
��?B"�_�_֤<�#[�.�Sɀ{�v��2߳Bf�5|��"�MA��sg2�l�pj3��L���ʑ�3/�z�B��i�����0<�~��;��U��#YG2� 	��"6���%�,�F��K)��@DO�2oPs6&$*N�r� QєSڟV �	�;y�xyǞ:B��:��Q1$~qZ��7�M��*�E=89�	�k�*��t���$D}�eLE�Ê����=�ԉ���A�_����O�vg���N<I,����UCy���X.�oE:Ֆcϕ���66�~��X��ؓ��֒�l .�g��h�Χf럎yo���'����{8l���M�0(�����؝�� �����,<��N���-�>M�`Ki�-K��{������7{�Rb��]����#Lh���'8���*���P�����-���e�7��s� ���~�r/�����홿��/���A�kVW�b�j��kW�IN��M����.���am��t����4�6�)X��9�M�9��^�T�b����c=�N������M-Lrt���e:��"�F����V�mq+�Q�w��ZLӮ�f�����<�O��0[#��ky �ǲ����ePC�3#������c�S�C�j�'�;"�K��՟�ߧ>�qz��g@�*���<��$��P���s}�#��7���ۄ<�LpRT�� ��� �HP�pL��#��2W;>���)��D�!OZ�;�lt��3�9�-��
^������˯I�8'ogM�$�N�h#�'���5�m�_S�v}���6�"Î#���
�����8	�G��;���$�6�����8���[<����נ,�X��&���bL�j���8�K����v��V�I?�����yǹ�5TI�[�l�2́}�ظ�����QE"���2��i���_ix||2�t=��-��|=[>������6��,��v�+1�����g�2ŇA��`u�P �����S�٥X����am$���/�ײ_2�.N���/F5i�e#
������G��iMb^���#���;���O���	����j�2��kLm��&]�XVB;�$)�)�SpڶJN�ڲX�ē��3��ñ�R�v5y���l���i/�s��_Tҿ|�v�X��h�K���v�rs�/��i3p�e��AV.	ƞ�[o��K:�r'�)3�����keZ�
�k����?�K�yV�6��V߾<8��\#��8Ѐ�Z�d�՝���v��*Ȭ*I?�c̍�Wq0h
e�jV�'�qf�8gl�F[Z��ڕ��jH�~R��j%Ƌ�a�oh��Ş^x�2�_5;��#+I]\e��	܇������"YY� C8[�K���A��Ɵ�x����VyT�(Yv��Ȕ+
{�ST?�:��7�Fڋs��rv�"�x�ݠ�q�P;���I�h��S��Ga�>D&A^+�t�l��E�+.,��\9;����zR �o���th���X"��t�h�>D��A�l�/V
��Q���<�R �\��Ua��ƻ
H����ۜ�M�lޓ	��x��j�*g1Bh+ǚb:��-���5��t=X`�� ��������N�=�J�j��/F'���e�Ŏl��� uZА�1�ˉ��h;՗h����J�JQ՝O�I �'��!\3$���LqC?߰臻�ż&��T��"C���9S�8������Ml�Z�v%���Ē�bu�T}E\�����6�g8����N���|����� Q i� 5ԺP�{���I������_�<�y�mc�*d���y ���O���a{�E,A�@S�z(
s��Q-ӎv'HْO���=vN�5�g�*���B��-�ږ5){�*��\럇��r�>�m%�?�3^���Br����	\����d�� {���p�Y�!���y)��_�����7�Fޫ�T��&�z{ñn�a�}��CH�B>E��he�_�+;�g�w�`��M���r���!7��4+��7�YWC��������~L'm���\�s2�צ� ��G�e�큷's��	���.)@ajST���Ã��Ak^��Z���Q4�:��P����FOfvSS�J5" �#�;>Ҙ��vt�#y#���K�X��&y����!�W�����9��[��'�*�M-�^�ZH�ΛTϤ'�����~������+�o�9jG��r"Z�a68��>�^�T�L3��8d���z���&֘�" ��C���L�A��:i:92�?�~#H�~�@.�aY�w*=��������'!�Z�A��9���E 	���a/�Ar���%�Ta�=r��j����UQpoG��;��ĥ.�'��(����8H�W|�g�%�qo�w�	�z�`���xk���I��{C�0��3����W
7�2~_��6�~�t'@`ѧMO	�L��e������%�-'8:[�Wx�������f�~���(�x�J~�iEd_˵����hK����|~��V��P8~��9�oT�*���������|Qb�ێϩ&�C+W�Kk(�\�m��b&щ��Ya�Z��[E*�I���S t�T��^���۶l��I�<�/�ĸ0���G,�/��Fh��h�MF7�����2'X-q�}���a�r<�hL�I����z���n^^Ѱl��D㠈�@g���9����y��ۂ�`���rPu�*����`m�F�@^V|�Z��x�%������gΚ	�*LW{�~<I�E�]��
t�C�+�T�=`��	RհC�w���m���P����/cH���kORe�v������r��"�aP�봡�Z��u��ʴ{G�)ӗ^H�)�׍�y:g�5�=�>�!��;��YʮK�@@�]�7l>�Ud�L�t:�,�K%q��,&R<kXf��*W���m���t(�:�D�iX���N�aҜ��gf\j���إ�X{��>���H����DQJ�>��9c�
��j[(=��<a�{#�۔�kv7 ��y,n+�����o����[�-��z.��Ý��s��2^�i;h�@�E�pg7`�|�G~N3����|�$-�H��/y/{9@����ɰ�Ko�k��f�J?C_����Z5�j�������;��p�+^3ί���w�%�?�Z��~���L�a��2�N����i��P�g�G�5���N�k� �K�G����ˉw���x�~,���-�_zk���e���s��_`��Cj�4�#r����u3zK��~�<���a��z�v��Y̢	��m�ٹ��2����n8�@Iz��A���i8�*0��P����	�z8���+A�,�=e#� 6 `�Y��)�l��đN�~��}����� �����YZ���K�t'����K�T1t���S�y��N�Ȉ9� B��m����g<z����cS?(��i�����.�{�UO4'�m������}u HA���Xj)������1��4������<�ߦ�U�bѧgI$ 
���`�
�&J*���V�h�o-�DAKlc��a�<�F0�9.<\���o����x=9�{:��5ƒ7�}��]����	�\��{���/�����f�3)�XZ�e���F��+5�H@+Ô�\�P���Bv���qh^��]�r��c��߹�g�Y��	�n�E��bRzvd+p�Ec1��cSŹ�׸^w����Xhbc�K@ܑ����M�n���Wx��9T��I�bѱ>��Xѥ�3�6�A'X%�t%��(>�|�J�/k�[��욚��W�%�D��P����s��nR����V,7:J��^b(��s��,�7ow���=<K��P�V��,z�7�6v�,��rH0d�B��3��x��굂�,ŲJ�%��6x��Cq?�4r Q�U���F ��ǯs�H�˯}���z|m ��όH�b�su��p��ě��L���Dibbj:�9����Hz�SO��u��P�Iǃ�)M��,�h��^��p(!N2��T0�mc�#(󮅬_z��nQ{F2��T=A6�ZN�؈��	#N�,�O�{�Œ��v�+��
g�<gx�vQ"�V�����4+���n<�À��Q���	�/Z��[���_��i�#��m�5&��3��e�� ^�GF�P�mO!�DM	���B岆zU��J[������xܝ@D(픲Y�#���aS����"�*��|�Ļ.�J��#C�i��� �^���t��b�{�ε;JW�|��eEG1��9�}��.��L2��
ݲ��#{���j�v�f�ft�ҍ�̟�*p2JS�����o���^+mv�U㏰�ɀnL����	dJGC����l� �Y�p_�D���$��D�FN�s��w(k%L���t:�?H���j8��sQ��N�OϾd����ᔶ������'��CPB�h��N�c���ˢ���0���CA�3�ƍ3��0�]�F�Bɰg�P�͖h;Fqw8�D�)��|v�����:f=Z�a��	&���>��O��X��j,#�}#R��zHrzC�9�5�U�u2�a��fl��t�#�%ެ�i����xՁ����`��e>.�YrԄ��W�=�f:h^��q�Bą���a�*@P-�3A,6��єp"+�O
WhL�X����hc��_�j���?�@K��]����C���'%���F�2jb\[C�%��_����&�a��m&��M�d2;����Q���D[��w�޻+w+������X��!>���͔3�E4�����%pH��G�#ie�N?8�\9�Xy�+�|)3G����< ��Ŕƍ����B$D��*h&9,��m�)��Y���$o�-O�����'&6��ʵ1�u�V�P�+?T�m3�����z���Q�-Vg�cd����eIC\e������h����R����RjQC�W�IZ%wZ8
�6Ӹ�)�Ahe���:\���	��^�k�k��@���&�}K;"�g\�s=���}-��<9�錔Z�Tٓ��'�,蔳E��g�7i�0P*����[�$=`Ѹ�"޽�?{��������2A~��	j��O5S���g��,����r��f��M�2�qn&�s�&�\�w�9ˬ8x]oIpRǻ��>g��F"4S��t�]oZ�K��>����|���}�'�I�.�]���&�N���Z��͔���Fq݋pG�x�O�F�x��g|���	���s�[M(E�e�c��:�@b�E;�v4iF�.Q��������$E-t��]�o	�(��֥Jf��R�*�`�Fs�Tҥ�_��n�|�V�� k�j�\�*ܤ'4����g��i�KArte�[,7W"|��.]� N��G�C���<@��\�|.,��_U�Y�����/�\q�{1�uƎ+fPi���$�#Ō�'"@S+y &"(Bm�F��I6)9���t�F�^2�>�������s�6.s����(��1T��5���7��\���O��~���*%��Ӄq�� W��*C�8��SB���C���C�/OI"w8�R�Ֆb�Q��Ʋ U���}iٗ7�*�
�Z'��>X<D��<� BϮ��z��vt�h����H▙�� �V,�"{D���,7 ��l*r���:D�k�q�#�����0Ygz�U.�ISA��Lֆ����y��_Zd%���L�;I��Z���e�X�2���?9K�.$��nm�N�ï[Z�����A\���m�������l�_�����0����}�!SXn��9$��*�2�����k!g
�p.lȰ�y��N�,WL7�u>���`��-R��GS�'� �%T��(�$�q�@�&� V�f�3�y|B��%�s�Q�8�D�� ��B�p�3�ht�X�|C��<�����j���C��V�agݻ�C�|e휕�1BDtɉju�j�����
y��������-��c�]<�Q�.4��B����Gd��#�B��T�6�c1Z�:�f�
��4E�L��E#L��B˗d����;W�:'�O�&���_�v��jj#����A�c�v���Q���5�3�Nl]�SL��s\��D��d8���2D������Khg�K��}��FL�h�6n�f
���h
��$��LGu�?-�$���<ho�rl>�僗5�?DZ"KX���8[�X�˲
ԡc�MД�ϧ[�O){�i� �?
�r�Z����u�f�@m�\�����0V<�B<�x+CJF����o3-9;��(gO�'�������n%O�9_���ք9\���Ǝ�Gw`�<�_�N�4�eL����nN��A��!�N���]�ڧLo�e��p�+U_Q�sG�_
/��'�»��e�3�5�Y�K��V�l7�B�	`�ڢ��{��7�
A��tXӛNe���ah��ۄhs?G�~�lu��W���59��ޞj�y��k�E�&��٬������0?ݴg�sC8G������I��x��Q�ګ��/jI�ge���Z��3a� �����}�x��;d�@�5嫋1�˙�X�M���v����YQ|����'Q����]~����jm,34#��0�7��)v������\\0#[��{�_8�'�H�*�t޹�{�����E����g�#j�]2����ya�w(>i�&�SX�B՝S���fK�1P�+\���:[�õ؀MV��	+�*(F�Y+��F�W
GګD��,���	6�u�+�zt
<1J+������/W�����ϗI�����Ji��,sU����/
�Z�VXS��r��D�]wp�������c ��5#����R��7�q��.[�=����bt��8��<D������G3C����(S��B4�I��g2�,iE��ٞ�m�Gdӕ��
t�^�Y����y����e�Ƨ͉�;��ʟ*s�2s��1�������2�7��0S��є�YpU�zTt��Py��\iÛz]���/����Rd�6sZt��B��q�͉@�py�m=���o����`{�'��6���H��C�L9�1<���cӶܮ<0�t�,�wۛ{���ñr�k���ї����&�ʶ�g�!���fxCW���1��X\�|�5C�*�Ç���.�\��o��j��Xҥ��;���g���u�2"Q\��6&U95 �2�o�� �*���ѕg�ا��/Y7q�m޽Q��#���9g�e8�KR{z�c\�(������Y�L��g^��qV��S�r�A��5}��
)o�W��L	�O�%�E�T7��`Q�4��K;�e�r��q^��*�w�5�F]�o=ᑻ٢�Y�+��~H�%�$���Ae5r�l�&�j�l|�"jF���jі���&p݇ҍ��H��г+Y^(�5�v9"���r��Y��g}�v�c�N�	�"�L�	�Ɍ���)]4�35���A?�#�PK^B�Y�H��}�Dd��Ǒ�`���t�7�i�h��$�]�@9ۗ��=--���[���4Ig��f��v,�=I8E�"��{;�{��c=A��$�Wb���-{�/j���}��F���͑��0�u�����H�)8Ր�B�O)qa,N�$��}p��Q7$��-�" ��U�Ͳ��5�c��oy:�̠U��d�p�R�p��Xk�I����9��p^���������m�i��F��+�6�j�;W5�Jj@��Ǹ���M]�ۡ�LK��f$¿SA���M3��~g��a�,���۩�r�~�ō�^��e�C��]��9f�|֟�!{E��8^�LO@�ׁ������p5�m��2��(P�rB' ��%��ׄA��>/7Ez�V�N~�E=G����q��J3�ʡ�$#�])$�w�������c��&,��.�y8�L�E��[4�չZ^LG�aoґ�4M(O%����j�ma�E;D�;�q
ɽ(�@,�����q�Z+~��;�M�MN�aX�0��X0��S�XR���%#e�X��[_>�7�cM��mi�����WՎaH�~-���kV�ծ�c��۠�ˢ܀��+ノo�-��=A�%5�?>��I����2�̓eO��� ����ߥ��jG�b�����ܽ���4,+��3��r&�ܗ/���z�:T�B
�J��c�e�_�!R+XMA�8��=
=���%�pG��́h��H)殟�c�Z���!P�5;�Qt�s�>��X�>uN(�U�w7�~Yhz]��<§����G����T빓"�m1�����Nl���y<���m����\BS�Y!���Y?����u��-��s []#]D�i��@S�ӫV�x�*3b�"=}���B6%.�׉A݄���<��9�T��Y���fǷ��DG���Eg��� Q��F��vM�+-mHG���r��ԥ��Zo��`Lq��L�u	��*��2N�汤�BҠMe���n�Wqk2A�V�y�Z_),ȩ��x>���"�Tq����(��p��%C뜼CWNo|�jvl���%`�\���a9�>cf���7V���n��� 'a��{�+q�p$���;P=���v��1���q�����*'�6���!�um?�(,/�����׀bj&O��"�� �(�"V	�|Q��ۈ�h���Y�S3�ř����%Lp:�tϋ*m/Z8'�Л�J*g�y��E���֢�����7.�*�'�r�3��������Q<7Y"�F �F+���DV�6?S+��Md!x�(A��=�I笓�{9�E�]�/8N��.��΃?�×hѣ;��A�;�}�q�������g�ES��\g��,��.�_v�_�9�9vkVJH7j!�)Ws�p��pu��j�7SHy#7bT��?��b,�/3�$t;�L����Rn$kQd�N��/p��)�W2N�y2���r^s�f6p0�����
>���*�������R?���!�{�ݦQ�����^5C'�	|m��t��)]�]JDI�u.�8�W4ĚY2���(�.�ծ�-�Xx�[�/c�>)䟸q}0��i����B�e_���S��-�*��)QB��m綠h1�|�y������=8���X�]�980m|�'�nPH	,���"ϰ�1�vEZ�`��;���:M����@�wK�yN�iv�]wږv��i�zr�ֺI�x�w>S��T A~�Em���iGF��W����=9�@{~�������5�}Ir�a�5��8��]���lB�F�8P�1\lI~,1�)Ջ+��Tj���6"����q^�
;#�2�ɶ+���R�A�4������6���	2��n)��y���OTa�`��*BG8x��:�B93vѫ����p,��K��$�4bG���(ir�N5���~���	�� ��jD���= �Єǽ�Y\�\7*�@��W�х`�ɿ�\��o,��ε�$���4{-<���u�|�tu[�I��D�u���l���\,ݾE|�������|���n���@���g�|��[����.ȸ�j1x'b�t�i�8���[����V�v��o���7����Ѿ6���{tWʹ���y��l����!���ة /\�K[�ܹe��͉y* �!����F���]�$J��ە~���C���4ۤ�(�m���V2�/!�{�����W�o�LJ��}�ĭ��	�kʨ��(Swڏ��-�d���_"�k�*9���ǋ�hX���b<��dhlg�OH��^�=�k�v�Byٰ����Ⱁ�`ߠw�&�w���o: dԥYs��8C�z^jc���;��n�HOd�ҷ?�/���W\h�nzy8{L��,�__���z���s�&�IE,͙�g��A��f���:�W=dq�娾�	4A�ϓ �g��RǮ.6V��"w�j)��A�-K'R%u ���&T�&�i��' JԤ���,6 �6�t&��ױ4��		���I��l8��d�݅���IcD�E�p���`%Z��,��H�v{��f0M�����1�Φu@�ZH�*u��܌�<1����=1I˯r� s�A�_'��o�Ŏ
ET�u#q���Ă�!d�N,J�7C!d�_G�Y�����Bv�
\žqY�a@6	�q2 Pyb&{��W��TG�ńJ�Q�����V��f���qE��d�>V	���W3���Il)�[����p�I�o�WR��Uͥ�����^�QwRx���U���$��g��ɞ9yꅩ�n�t��z��ɐ�oE����R�2�ȑ����b�K�^�Ghj��6yb>�Z��o~�<;��qd�k_17/ͅ1+��:����@R�AO����2N��Z�-�%���S-A��M��0���U#�Fa؏/��[��d��Z�/:1͊���sF<��O���Z*��ٗ�����h���f]@kF.����O]�G�5�_����$��k�C���P�j�G�|��.8�Z�l-M����w�t��UY.����]hm��x�]��t�kpC�\�c@�p?X�"߳5X(@���[��x�c3DTe&-��S�s\of-هA&���B'0�δ��au��]��,�2���)Q�j�k�W��:~��#���B�b5E�[$넴 �9�ˉ�|/l�Z���Y��.�6S��u�?CDJV����D��F�P�%�g���\��T������15&{���q���T��Y��1[R�}B����*�8)|�&���K�?
{��*y ܮ���b����3K����& �?у`%��3���'Q�R�"	�kPD<�	��\�	7���e��`�U��I��q�m��$҃�9�3�Թ8ʨH�#��5�ӢK����j~�Xw��K�m�}z��m�@�h�k��Fb�O�=��z��j���M�K�&U4�)�˲�Ø�����g]���oŪ�z��JLѽ��)�ːpR�z��e2�}k�
=�9V�h��*�etQt0��]
n�-�|іqc@~�W4����%��'�:�����v�
h�$.l(��I�U��KmF�^�_�2�� $7;����C���Z��`�4ͅ�)	�XI^+!ySy��clB=�.��f}hb�����LPE����uuǫ�=��]��M�L���^��NU���C��P�r{Z�>��s����)܎�L�qh�~���+�lhH�`_�	G��[B�W������U���:�H���ް� x֗��uC}(Refܷ�X)�������QpF�gH��|�����3��t����Vw4��)��=�0�]����Go=��0+�؝���v����u����J���T2��� 6����P�\y�B������FM���{,V������?����4��V��j�e�kPS�D׷�\���y�L�*��KT.'��-���L�	_��2��N���4�ַ�Hs+C����R�F/+/W� i���"�GrY�_MT�u���^j��z���rX�r<{|��7�Dߚc%��E3��m&h�. ��e����I��T2_�7�B�0�?/z�:~8��j�Ȑ>P �{�ѐ��W�M���H���ҡ�O����Y]�ί�?`�ߞ��Q7��.��7��e��Ж3m]�3!x��i�� ���e�Ro�>jKi�er<K�;��;X���@!�b}c�x��	�e��x2_�GՆX^�P.t��N�O{aL��h���ۘu���Y�e�1���4�;�Y��)���K�綘{���N�<G&+>�ת�b�9���+�.���L��CP,X>v�B��rB���ު��֯ ��X=�/z��d�zQ�wB���\��s���A��+��S��r�՘�\$�:���Gd�G������~wƅw��NQ��I:�C���f��gᰨ��D~W��[6������ܔ�b��>�/��=߿����ֲȵ:����k'�/�xh;"x�$*�|�U�V�I֬%{n[�$�{2ƛUE�����G�s�K@���0Z�~D���"�w�꽽�x|i~2�3DL���s���I#S5�L�40��Oa�w���.�Pg
�N��{*{c��8	�z�1���@ަ��.�"�ͭ�:�g#���S�1��}.�A�-���&1 V�ᖌPj9�=S!��c�0J˝��8����O��	eg����|+�z{F�f��m���P��)�/��{��� ���!X��h��hx̱�M�WRd��t1�����rXV:��Q�#1��-��B��Ԭ�BI��@T�h����L��{�u�����V��.�c[�Fs:�i�
u��u�d)ʕ����j���'�[~.��_wP�i����mr�\W�$^��{��jΓF�[{kb�IRRc+_�$�LM˳�s��?=��WJ.��h��q�i�v �K����Q���~�"�4�
銚>����r�ag�P�%�߯e��9,B9�ws6��0�BPB��B��M]WV#����8'q2����cO	0��.b~�[ْq����8m�]��.r7�������
�Q��vi�
5"b=�l�W�%&�$5n��_��7^K楘O�Lr�#_z8 �QB�8�, �dU�k�rO�'�d3.7���\P�� zJv����9 ��,������� `r�W ɣC���.A�	���f)�x�fq�:����v�k�oK-+�����@0�pk�-��'+�M��j�(�ǎ�^�������>�Y�7DQ�\�����Cjg�=��)�r����T�䔸bY^[��EX�Tի��)�&��A�@�ĉ��7�C�&k�*��\���]�_t�Y/���XJ�P��lS'�L��q�{V��^3�3�$�6�ņ09o8z�����C��TI$^�h��?:��Ry�����J�� ��VB6�����$밼~=λ)�q�䬨}_���.7�.sŚ?ˁ9���1�0V5������ٍd�;�aD(G��6�m@Ň4��~�DX��V�Y�)��;5H��/ץ��'ܝ�k�W��x�oC�b H5�]�կ3�<��t�K! o�s��&nH��o[����mL&��ns���!>�LM6����LZ�F*��%brj�n.ĺ�R��|�?@s��w���<Xh&���
4�X<|��g`��-IP����+0�	F�����SOH����R�AA���.r�\��c�}A�x(bF`v�fI;5u��Y���>4���X��`H�X����Es�O�3Q:wF�C6uV�}(Nȡ<�$��h����`�e�s�cf���x���SyF�ټ�S���F�+܁��Gα��ʘl���K6��ぶ�I�{�+(q �Z%��8,��E��o2H���[�Y!�F%6��[52�����~Z���}���Tik9u&g.^vt��C^��i��%�?�����==���諦2ߑ�{i�25;6%N�s�'3��A4�p��U%7�#g�F�n�`�X���{���T( zt�P[g��Ryj:,Be�M�N��䰷{٣�h��0��f3��y���M�9]������$4���T���ˌ��LI�5�����9�SD�TU��eYO����im;x�9v�B�	�V��~[�'2���fd�zdt��0�9s���>&��;)��6�pT��<�B1Î�g1��b<Q7?�ʠ��g�u��E��(f���N�7*/M%�kN�$}�*lo��X��ϞN?�;�Y�m4;2�<
"�I�Kmn}T�"��0*��y�h��a/�͖`ݚ�-����c��5
���^�h��dv緛d�u<� �.d�uI�[KJ�Qe7{"�k������p�/�����Kn��>�����Z3�D"Gf�\�����?���8�-�כT�PF�9�1s��%m/��_}����U�ŀ�z
N=j�[I_��aJ3�,�I%��8�å���Ǥ�1�N
�&B�6�4:�"��n1���M���Ge�]��j���z챃�ԞnW
tS�B����t���	$�@3��b���㪶u�A2gr%̿W�Ȉn��N�x�?��'F#�y��c�[Pٳ��·dWU�m�����'	��J(CC���]OϮ�b���Eʴ�>�6�:NR� D� �kZI�|R���KI�L='L�r�1�K�/R�3P��X������pL�V��(�����u)`P�����hI �[Lb��o�̉�����;uJ��4tK��hV��9<U��=hg�^�FJ�l\��S���nQ�nf��PJ�}���6���O�d�`�, ���R�HygQ�iq��u�끄��}��b�g�k	��AFo���?p�����y�U�v� Q3~�Q�E [��g�Iun�z� ,Qv�!f�Z���K��gC��{Q���t�",�4�����:O���(.��B�1� q[�'ckM*�`���	�7'���U�`�h.{A�Tr�T�N���n6{T��3�*1��i��\)Ra���A[ h&���ɟO�lc��g{����k�JkK�@��^�&���GNFX`�AOp��:+�Q�I��I�b�<3�e7�S�5.eɯ�Q��c�A{����|���Ns|Y%��������i3$LL4���cv\$���V;9)$�T��G3w��6^�D����H�g_���?���2f�L�{;x+,;����sNਚ)ύ�0m6>xYi;{���9� 튉�������i�9� #y3����P�Wd�qm�[�+!�)#(ǖ�s�������M��Էb1���<��~t.�n�@L"�u����N`׎{��ՙݷ��B�}�����lޏ�+й,�>)�d`MShS���h�� \	郕=���P���LJ��h�O1J_�\'�l���~�ԆU�7ڈ���V�m���k�T8�r:��Ș*G�����>�a�!�TbUȸx����X1�i��1�#�{���lA���&����r�F\M�f�68�S� `��<r��#;����%3M���壞`T�8�{�o�W��^\Re��vL�`4��E�)1c���2�HD��L#Y�n�(�ׇ�EW��|eU�d�Nd��ݸ�����x)n�I�U�� ��S�JB!i��BPI����RkHӾ�
��e��`v{�?�Iq6����'�����K��%�
��4I�m74�̞Q@�PY�~�B��A�2w��LD\Ee2N�x]�ơ�0"s�;��5��oa7��� ~�E��x�@�d��,�3ÂE�������*/�"8$SF2-b#��u�Igk7!<W�'�sF߉�2d��ƭ[�`����1��sa"����ٮ�Q����8a��5IT��P`ר�G�v���
��1�Z��7�Ct�3�9��먘^��2j�]���h�^�_EL�+Ѷ��%��^��� o;M�ӏ�CU�!2�� �`��:�����8CC�ʣ�Qy!#�y��8q�6t�]����/��u���N@F�Z-(�C�o�o���]�I��
��0��zzӎc>����d�W��@�����4ە�s&�h�嶄%H">~j廣���!�Vw���Fu��ab��#�9d߁y��Q �M�a�<��-��?q�7���Xk���K��RGD�U������1�J>�e{����<�8���MK�W�ҋ� ���i��6��'k��VT�P��a���S��]Q8�v�ٕ��깵Z�S蔌�HlY�QA�r��`�j����*�v0b��BZ���"���5� L�j[�\Y���a���E_��5��̹��N����/OR��jiq��o~|a޾�߶P�������
3���b��J�ؓ��VdxZ; Ҭ*cO.��D	�̾i�����/��Z��v��I�L�+p�Rڱ�YI�a@�����B���H�jN�k�	i0 ���~t�m�373_8�0'^�����k�M9�"�6��X��l#�gz��
�����/�x���yLm��3q���<���tC��6O0�bf��kb��:���ҹ5�G7A_dn	���f�e���l,�y�	�9zU�ɲx�<�����e�D�Ϸ{^V���?���
Y�
\ �����A
�em�#�]�~��;�]J	�F��ɵ�-縻�K"a5��3V�"栵��|8��fn��ธ�9�1��u�/����`+�s��Ǻ��Tڶ���>cD�^L�x<�\�Mu1����k�|�����;A0�؞��5�W4h�J<�J�#�ɋ^Q`6z=�С�i�j�h;nߨ���ި{��0X]#q�#��*�FMMm�~��3"y��	=R�?T��:�G@
������ⶴ�R.!���aO��y�[�|�h���^aZvj#���<�Ұ�;�R�:���� �N -7��xD�5��Ӯ���Ђ1��K��d�Gӡ:T�B9uwhfyY��Q�e�)7�W*�c�Úf��S$u�{0����ŋԿ��g�G���	��߹H][@�@d��͆]����lࠀ�Q�O�,0m�P9�N��O�������VM�����'t���A)p[=�BZ�����]ch}� �W(}4o�y��Y�@Ep�R��xG�:�d����P����i������$���d�r �2_Q�ן���=�5,[����z��xA
����� Yc���Hܷ��M,��~��Cl3X�if��[�RѠ֔V����Z[��;l2�$��A�?���כ6��1\%�o�Lg%�;�bs?M�V�z�J��8�	M�Ƚ����q{u~1W��2�/>ˮ�)e�\��(��-��A^=�"����S��`���jP8�NMl17@�~�Ç!�O}�m�?@{��]s�7<�Zd�[����\��y���LKCq-4QY4" ���E��X�.2?/��͹������5��p	���'qh�F|��M�3��'= ���,�c?�@UI��%�?�����$J�B�7�R�M��xR�S_-P�Y:kO�A ���pT���ǜ0zF	���B�3g�� �$�iI��T;��*���j�3����3PO�!���RÉ�I��a��R7�n#��)���B �w���m�Kq i����N{�n���\?��p�Y�fY@�8ﭾ�gѺm�c�+�?%X6%n�z���t>&-5 �#.����!\����ު-��ua��,�õI��\Pn¸�㼼�r�Zp0��A�c�`�����&��������g`��/Y7����"^��������ѣ�%��)W.�c���Uf��U�*�q�ٔf-�V0u Dp�Áv{	�OY�2��t�A��$ ���ז����������>�h���>U�ll���h�BO3 4a�xB ����/���b-�W5I�� Ԩ9��g�Nu�q��zG��˺��)"�t�����S�Y�jQQ�u���ԷPo��U�T�����ݶ0�'1%3GW��蛋��%"8�}�W�/��k�<�Gd�Xʑz�}�}��µ��'Q���&ĸ��-��ܝ�Sv~�1�$����~���'i8"�b���$�=m�|��E����]Bt���a������[2�d��k�٥�r�Cڠe��a8B�A��'em�����!v��!̦S�t�`�2�+�Oh�x�1��UYM��t�Q�r|g^�15!ί2��ʃ�4����D�_���vH�@��`�;
]��m�#;UB������~���y-\�{|�Q�v̂�ثi�.q�Ɉ��-7�Go�w�W�f5x����1�q7��O�ߔ��y����<�n���Vt�?H->�2���B�E�ȣ�k��,�����g�+�h|�[G�d���}��|B�j��=#
7�ܻ��6[�e�����4��;w�}e��B�b��B�8���t+��1�0M%&�z=eT�2�I{���F�+Wa��n�K��v�c7�G�~��:ڷHUL�j)���V̓_��$\�_�&�ufW�/I�u�.w������i<�B-��I\��sԍ5d;T�l�8�U��⽬c�1�M�Jwg��A�6Q� =���N_��]��l�'�12A�����!.є�b��Ȥ,/�d�f�c����H���϶����������1�D�
t�@K��:Q�D��L@�]vb�^i����2��D�Tq
L���X!�7�AY���jk�r��M���b]�<���Zp ����5}@6slg�:(�}�]�̓����z���;�Y#d�/�X�W1рS�f<!��cɃ��d��b�r�d�!�`�t��`"^�AC��` �O��·H��l��6E�-O@��rW�R�O� M�$/�F9���^ŗe/���[��C+��]"�ʘ7Y���ieH�>�W��gx��$'�����8l_!�$V���h�\6�Lv�.�u�h��Q�����<�DM�ɸ�|.Z��U3�9�72�E! ���rd�iZ�-�F53b��'
<@	Df���j�=&P�Dҵ�x �>�J�z
΍�4v�7�����v\��T	�j���Ub?�^�G�E�~�^y�b��m��gsYF��,�1&��u�t���JS�͘z;S�,�x����ǲ:~u�?�(�r��E��u:�9K�	J�Kw��tA�b�Y�qf���ؼ�a6N�����ً	�j]+�Rm����s[�U�甤���� tn򂻙C�GRTf�y8W�˔����#3;�g��4!���į�w>Ƙ`p���$��򇰒�:9j�dY�N�(Ewhfâ:t��t��� ��ż�d5�ɀ��l���s����..��Vю����D>r�^4�ꎌ1�8�Ըz��9'R/��;��P����/.�'��5@�3��ٞߩ���x��	������LyՏ��{��f�<a�y�D��p4kD��t��O51���i�@=�/�p�(><�'��2��}�����ݛmXPW�Z�O���f��e�ѣ0����xh�XU��|
�_�k�5n��i�&q���w�u��J���8Q2��$�^�-��z.tC+��A�	ċ�u�"����b�54x$��C�q���l�l�W��rV�R�,��DO��q	Pi ���g�^��M)EY�}!����0�_Я�@u3�U�r�!�-g; =�p�Vح?�S���;�b�y��(:����#$���)�[���?��F���aU�S�L���<!V���O�©^��*�h0������H��
�w�*_#�7����u�!9W�}�lFý �t_k�	�����Lqb�~el2�(H]�bT�W�I�r̙�ȫΦ�d���Q!�,�x��ŕ?:¥�rJ9�TPh�ۇ:I��|+���"��@�)G�Z����PmQ��Xv��;Ky��v�a�$��T��(@a#Ӿ�J}:�&�p�&9���;x_�6��7|�@�ۆyB=��\���SLTá�׷���f��j�����O�W���^g�c)�B�D*F�OFRi����$J�LŕE�G���&����P�oQ��{MȼGB�Z��
�2��������D��R�F;�mHʴ��J7Q�e�F٫�#�3������>M�����s��/0�v�eB4��zr�t<��F�A���?x)��Eu�w!���*!2�Y$���5����^�5I�ܘ����T���zim�3F��X�������V {��\�L[�P�w��i��2ɳ����;k��Fs�X���)�O�c��6��5J�O!��	#�7��7�u�����{���F=\`�hX����יBHv�Y8���{��oA��P/9� �W�8Bp*l@����?�̑C�� 1+��	�B�JʌcvI����K+Rs7��
#�Wｖ�Ld�>7���Ző�3-!a�(��A���ɸ�q�fc?�M�,�����e-��2/�a{v����(X�t��!�&�*S�[��D����͝�O�z�$ra�bĴr�6�>��.Εz��u"�p���J��9�yB"��$��(�����wl����:�l��
�Ԩ�������g�E�����3�[� {EЁ�o�����ӠnCVzS����ܫT�EΏc�5�ms�g�N���N_h눤��Y���^O�������m� N�XKS����s�N�&��C#c������;Y�l�ihFR �y��	:��w���|�ȇ��$�y��4	da����t���ϰ�e�s5����WD�<n�&!:I�m��ea�����?��"�	���LO�^c��~b�����ք�[MEk?�^��
TT��X��To-6U5�8K��Ř��pR���,��l^W���%4���g�G-�ާ����+�w�A��Z�p8ۈ���GV4�?����u��-�`#�щ�p��Q�E4)o�o,���։�|�V}��Q�!L�����B��J@�?��(���O��v޽��<ۋ_���}��R|C�KUa~!+�>J��l0֞p�'� �T�K�*�e!N���ӄc�UbWޟ��~��6�u���!�=���x�`$�]�'�*X��7��Ԝ���������H��P�[E�h�<Q�w��G(x��v�N����_@x�Qcc�\3������	u�;X��k:lF�k����vhj�&����t�3m�r;���v.�����{g�{Xt�
~��Y	Ι�YR%eQ5.8���*���#�Im���,Nˏ:��qq*{��K+U������_.�Jޏ%�&4�&_G�ފ���@�3�p�8�Y����a�|#�Ŀ4x7q���a�riqF9�+���A�U��R&�P�:���*�2O��"����0����=��J���9q0�7�v�F��0ye��#x�w��S��	j9��k��Q���ȦM*:R�?U�3�N������A��b��^k��-�F�u��I%"�M��$�JV��W���]�f����ی%+c��n������J�h3*�s@���6dy�d`}���@�)Pu�޻p]$�`��JA��$��p�'d�!al������!��uh,��\�-#;&i���覑MbE`���m�X�fЊ��zi5�n�h��ODX���^����M}�H�R8�-�F����Z�/>���!g�L��D����pHz\sƌ�P�b�>C�YjQ�������^��H�8��Ʉ��Aq۪����Z���ڶZ�f�P��h�E*Y�DZw�Ԅ$�����7y��ŗ�B����@�?ʾE��Wm/C���T�bk"V�`n���X��G,�&=�$Ԡ�@��A݄��!�r���C��}��ċ���T�����-�(wmf���~��W�	�X���z��>�,���Mt�ͯ��g��*:��I7�́��E�w;�i`�KaJ�Εԝ_�h��k0[1 	{��X�e��Y&Լ�u��m�'�	o�*9uۭ��P[���#`Kq7���v�4U �.��u+t#����tMʹ�`j�,c����4��z��T=c�*L��Y+�M���r�ҬP��+S