��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)�2������2p|�t��-�rd���8��u/!���l/��ɲ����%^%zMݎnM+��cX5Y�<RH�ʹТ3��1U��Q�B��{o|�/��W�:*�V�D�A�e�����D\f�%��ז��j�p7A�c�N់^�]u��Uږ�dK,,��n*,�O�aS����D�0�S%�=�X���Ljg6c3��~;�AV>���)�L��⍙4 &i]F,� ��<"��duǝ��W������ѩ���Z?c�t�� �vS5���(�KH=�&�GSkS�/�"�^خ�u�ߋ��q(`Ǜ�3���(�#�ѮkR��툌(X����y��=�Ԏ=��`�OE�����a.o���o�O�����~�$X��%���2�p*r��ap<�	K/A���g��Ζ|7�4�qR�	���4Ov��.����\�7o~�m*�؂�$[|r��i���|����a��Z�"�k��ՖQ0/9�y'���4�y�� ����蟉Dz|��5=7DX7�kĦ�~Vآ���Rm��WΫ�˓)z+:���d~V5~r%E�����V�w�?g^q	���c>job� ��5̰�h����$��s�Ը��0�J�d\-�*��EqgV���V�c�幩/����b�U	@Z6�]U;E1D(���4��{[ [^p�4Vƞ�'�㫸�M�
�B�2�vr��r����
��^��yv�QNe�ƏL�uK��03��ƲTp�uPnP�bT�<ֿ
�����ރ�Ē��u�ѐaC�b]���ݪ��P��qxdc���kVa��t��G,�.��DJ��j�h�¥Z({���$z�ln��G̜��,Tٟ,׹�j�v2v�N���b�����k�=�>�Zb�YU#����:h�c)gqW#Z��z�$�:����/z�y���<N�v4l���x�Q�\�֤�X����#�#�?)kS|s�g����Ֆ�WU�w��J��a����#ȯ[�W�<���<c��Q�"���P;�i��z�x�� 0��n��ѥ�4�9_���b_M��`>Y�Z-(��[;&B���*�O"b+�飍�_(����B�+֭Wy��ml����mD�~ղ��>JK�?w(��b{�G���_�G]d%���>;cl���E;�N�.J6�q9�4
�!����0A��6����XF<@N>�饖�2���A��\Y�A@�,�W�j���&z���*��Vi%�-פ<Wї�z�qf�+���q��i��p5O��O�(t֌���/�/(>,��T;8�Û���Φ�!�]$�lu����{���G��%��l�O�z� @z��Ɂ6Qv��'Q|�6�}�d*��>eg�_�(�����Ls;�'�M��^����_�*��9H���߬�e��D�T�L�OA�?{����
44B1=01&�d������L(J��\kc��SL���95�Sv�_I
6���M=��Γ;�W�������ЉBTK����-��zѮF�����$�8:���S���;]�f}{T�4�-S$a�?ůSo�/!�i4�W�>#`���62{�uW� �N0����R#��B�^�BOL��4��&��[����jU��/�aDG���h����Z��u���!���R�E������;��U�wcF��
V�|R�j�H��ʥ]u�5�0U���d?2fְ�q�8����������+e�wfO�kC�S����(���Rt��j�Ή�Iju���_��h�΢���v��.������Y��(=��=ᖄ�l��z\-����˴�	q�
q��1�R�o%�/��r��H�3�}6 LKK�+""��QMonlXk��Z�%c2K����͞@Gzp��{�&�Vu:�8�\��H�2	C#�,����K8����cm��
Oo#����F��n[�.:(�=��[��w����A|h8V+i�eJm��B������l�R��P9��%Ps!������*O�G��o�w��(��(��NJ3%�>R=�_uc<������Y>@DE<p�F�haU��W%�	)�>2;�Y��UՐϪ��Oq��&�EB|���~j6�(-���A5��Ѷ�ĨuR�S�@�m���O�� ����G�a%�K��P&��'�-5�~��"�J�T}X�x�o�2Z�U��^�V�>�4�n.ü̫���sp�,&��Q�_��Q�+�G��I�������\hG�!���m:�wN���3��Ɩ�����޾V�J�o��2�YX��g}���Y��kh�/t69����Ic�A�w�lߤ�.)��%m,�`�>��i�}�۲2!BG�|�z��[U�葉�1v�ﰭ�e��n?�l��#�ʒ����˭[h�jˎ���b����R"'\��)8ɿN���c��$�3�h!�/M��'���2@���U)�BE�D�M��l��:1F���@N�|�R�#<7��a�O�� ��rV���]]��r�eB%��<�$L ���qu�m{s,�^�c�9p�(AI����vUS�&�s�(�
��� �H@�S9h�%��Uq�*�^�f�2f�V��ھ���ݒjK�a\
���^���C�㾷����%��-�D�7sM��I�%����L�F� ����D�%)�!�(�̗�#@��e3m�b��\�.��w(%~u�6[��ws6���H������!�x:���?T52n�"�\W�ƫ"m�ǂ�o�La�%+�7��q�5���A�εC�Ĥ�,�+�P{���c8��)?�R�H@��{<(��d�8=U��?H���w�Q`
bCk��M�F��Uҷm_ �	��cٙ��D5��?��| ��!�}7E�'( Y6U`l��	DlNZ�Gpb�v�Ƽ�'����ѧ�&B��,?w1����`�� D~�k���?5�vrP����µQ)5��E@<�Шwώz�@��B�����*��l��ݒN��)�D�GH�Q	Y��^�5�|J"�l[x�ء�,��@��"�.����m��FT݃�=%�~�F65�����!V`�s�c�q Y�֜$�Bc[]`7�!��B��I�^�Q�P*%5ǋA��Z��s���!h���X"%��m+X�l҆~��f�D���'.��� M@��X�\7�~�P��Zu��2�7��x)I�ʏy��D�uD�KT*�lu�*��"y"0�H%�����8����g1Sbq�뷱�S�'�ȭoT���:U��\�_w�Ar��%zOa��@!+qt?BZ,��*����lGfGg�DָfTK�Du\�I�{���T!��;�"4���;G��A���.�m�};.��ܿ��%�x���M7�r7q�&���'�����@�\Љ��^8�o�D�OI`���3(�;|E�8���M�XZ��d�-ZX�Z8����J��b
�51��	�P�{nh�j������Z�3�����~��4�����o�kS�q��l��*�� �ϋG^>�!�g-�YJ�{R�T�xtF�ι������$��#۴`q�w�v���k"��K�����ˑ��=����d4��ǟR����Ϡ�� ĢԨXsW:��e�?�+��v�����B�~�7�~ y���j8���'N3�ê
���6b�~G>�<펊"w
�NR\F�����uڒ��z$|�
���)c?Z2���&�������F�]�>)��43X!<>�n	��c���Vz{��($ZV��=s�ￛ*�v��eV�	w/y��M]AgL �SH��1Q�hg� @@Y�A�B�.�}��w�L��/Xۚ�~>͉�އbb�H�
84
����T��M��6�b>p!f�����+\H1u��hY�S�����M�	%��|�?;����T���� ^�N:_	�M�����$��yK�`�4�Ė�N]���+A%g���->��"�mI9�)w�'��;N�#�r
�H�Y�4r��H��{jШsv��(���&S��%�oZź�����cֆ5�x�?21��3�@�����
�6�C�"%�(|����_d��P�}�D"�Ɓc.��1��TL��2FmV� w�!���@��X�r<�Dm��ύ� �A>�g�0ʴ���ۀ�?B\�f�7e��A��/
ZY���|.<<-3�89�1zfk��4F0��>3L�;�.���'�+-�m���j�aJq�T�j{�(��U�����i촺�'�0U|e#��*��E�nd��H	���M3��6&�G���� �]������qc�j@x���+E��)��tq�əTA����{VN��}��5).�{=m�ӝ�'[_��<�b�a�cX?�*كw�}X��?�ǟ��|v�:����W�ر:��5z�0*
�ԟj��~��A?��_ۗ��wX]j-. s��N��p��=��77@@�����
�&�g�jx��!��QەȻ�u�Ș#�,����zpRe:�LJ\�/KY֑k�)ד<�9�H���UVaf�x�,���{��rCa��N�Y�.T��_Q-�E�I{l��l"Q�]��E0x�S�_�����02��ȶ>qf{.Q7j]�����.B#�MTnm��c��}):�1�*��Ѣ�*�r&�P��,NЛJ����gC?y/9�`L��89ʷ+_�&�[�K�6�Rl��Ūt�5��B�~��H�No�n�d�X �ic��b܈�I���v.��dcF�e��ڔ���Y�B�,�ꔳ�Q�n�r�ɴ�2W�fvg~�-� td��z�z��f�D���E\����+�YIlse�P�7�ɒ��P H�+zak���mg>�s_��Q��-����*x�p_ij�E�}��0��tpƅs��b���@�����Z� ?��i{��+0w���r����k�X��8KX�)��FC��+V*�D
@C(a��N<�� z�M>C~V�[�s�u�By�s$��z�Fj?��X�Z��9Z�i����؞���E~��gDR��?���g��Rҥ��!1�UrG��4hr_ř���=�x2�� r�E	�*@Zb_�߫)�Yn�"���!��A�m��
 �����d�#m��ᬃ��iu�"��L�k�fX)��+��dp¨ݾ�KX�a���tmiq.�édo����=�7�'��h�"z$[#Gao�;�G�T0�N��m���F��A���g���}O�2�F��1���(��b�D��AP���L���Y{��'�.`����ۘ�?8I��n\����n�|	8�<G��9wf9�,�dn�'�.l�*)�����n_*Q�&o��K���m�����AnT �s��P���a�B�]3�F�0>�
�,n����]K^ӟ�bJ�c�yp�;�m\���Z��NM%ZQ��X�A�+XF$sn.�+�RK.4·�t�5��bw) �8SE�ZƳqSE�RX�a/�
�_MF�T�cgP	����p��`t�&N��~�g�T'�Q=�\��:�5Bܰ��G�
Ҿ���JyU�8���9g-� ����	fW��")g�#����s�Y�k����޼A�W����Yg��B1���-��-��w"�:0*~)ol���A߅�F[�"�x\e��������a&�$]�U��I0�^�<S��$D��8W����uwR��>�	�'�t�z�%�t~]�����VlZAb�����^��u%n'l�.�J�zAt��l�Oh(�|��0B3<s&��b-�ڷX���!#�WB�iV���2��U�C��g&i�P)�8+/�@�����8���肏9���}@�=�s[j���T5~Yq�RlY&<�'�U��BW>�I\�N�;�u����Ot�(�=�v+9�xӥ�ʙ�kg�@g��n�5�kN1��JA���v:m�@Ir`I�Xj�qc�10�I 2�3�+y����	�/k��⹄j�"?�*�����b>��Y󯰩�:�&TS�Ǉ��X�E��Pڲw������8�
h�Gq6�h��|Fp��Mu��цWW��H�+����H�o��� h�`��\vm�pp�����E��!H�H�L�"�D��U���8�;�iiP���n���z�"�[����@�Lz�LoF'���y:�.�׎�� ���������8�>P��ʑ�q���ʜ@����n����A���?��l&�ґ��)~ah��疽_Ώ�,;FA ܝ.X%�1v�T�Ӻ5�ym������z�`��w��=��;	�gb	E?�~]��0�:_.�u�/���$����n�ܔG�hi�ҙ��vזlȊ�O@d���U[�[�����?%�0݉9�+ѹ��B�İ|?=Q<�yg�0��\��ػW��f_����)�J����}��l���k�@G�A�����0/=���n��t|ۏL�{�Ea�A���%�Ub���ơmo��2���6��9IZ�|�r�����������!}��h�3�E5\�
�n+�F��*��U� ���9�y����40+ގE`���|��;}}���p��D�<Ę���S۰�g�J�	r4r�.޺����n�o
U��j>�%���	yD`¦�EwXTY�}ퟖ���9�Z+���q7��^���U:5��i�O����4�e�<jϧ�k!$�?C
db������ۘ�y��q][�.Lo.���j��a<A(n3tKbX�����,�D�?s�(4i��w�����:'�g4�K�e������/|�)b����3�������t�5k�w�p�7�D�C�ސK.7�I�����kL���V*�_���t��Z�(5�C[v^���	�S�)��
�d�$a nMv�2��Ί=��g2}?�_�J��dg�~�sٔ��;�V�������/�1k�)�I��|Dq*�K����P�؂J�0q~&2�q���P��[[�Йh@�ݐ7��.���O�B�dч�Tm˜���2�u��~�D�ګ�K2-IQ ��Uj��4�x-�f�.{��; �w��f��'�j--��u�vo��1����*�3�1��J�%F�t���>_���3�}�Md�RѨ��0J3����<��hE���in�����?O�7��C�\8�Jg10>�
��͹d��f��g��uĸ��;�t�1��	��P��^�o!r�_����{:�.5�˫�=O��m���S�X��iUf�i<�D�^��q�0��?�!�����]�������_��YNy��Z$&�yVb�
�χ3b�,U�a�����?2�}˄q����#��SX��G�w�Ϡ��Kn�� !&?9�O/�21 ��brv���~�C�:�_㴢��1a�6"?51��C�Q��W=�y��N)��;�͓�Q��n���(BFM����9^e�gH�=�:&��M�~�^c�8b��P!�ۥ��s>W�P�Y�3�z���ER�q��I�$B���u���!w6�I���(�^��@�M�w/�����v���h����E��˅[�x�:���2N�+I��K�P��r=_�p����m>̍v���?�>S���:S�aW�F1��t���i�'�[�g}┄�l�;N��9㶑sXxZ;ѫ�{��|�^S���um�އ���S����x�A��u�Ю��0�|��7���hw�@6X�� �_��)U����׼e�{S����x��H��q"-6ʫbg�p���l����<4��&|tT��UӒ:orv�������gd��+)��9h����w�Mp@Tn�:)�z�⥇���
ɺ��n��B��"��'{_�7�Q�KIx{��F�.,e���jp~�OԦ��)�䟺������*�{�+��U�������'��~n�HyҪJ�WMȉ�_$U�n�f�G-]���NO,+w���q����)�V�fQ��W~���8���׀V~ܕ��>��Ζ��@X�	���H��6�o^�%����C�v;��&�[��<�����p�:�9�Pj¸�� ��cOZ��R�����9�1BL�>�V�'���»�KQ\9$MoҪIy��߈`:�������p�[��f�}�Ar���)�կ$[V�!wp������+�Ŵ�<v�<r=���������yTa����RZ�
�,9�	/��ɚI���`�0	Uy�`F���M���˒�2>\�t�G���6�I[�.Ц�y��Kr5K߼��'����*\86�	.p'vV��)ͺ���!]6D�[(�Cm@YD6Bx=�hv�;�pl��Px@8�rI���qBN��#mDg��Z�}w�W���H�&9�\f�8���+�H*�v4h�/����:�`H���r��`�D��[9ߺ[��+� �-���h���UI�f��U��CcFx���#8��uV>b{��s�V�!�Dۚ����X4̫�
��׀+�<�JD0v�A�O�n ��&�9�cWd�<X� h���i���|!ڥ+G��U,�U-�d�[P���~�AkMg:���Z]��ZI�^� %�O�S�JvvuY�/B�BC#�~E���J�c����`JJ�}��C��F�x[ǭY ��@���l8�x�A��y�����*�!!2Bc�����;�WR�䤽����ˡԩ�W����^[�L ������f�'�_��Ƕ�;�g2/��A� ]KN �䞈��}�1��{�??��0�:�=�ˋ��=	��ݏt(���w��[��D��"���r]�k�k��-GA~5�j1�:�Xc��+�4��wtU�Cg�x�0lHE�2i�>V~�ş�����oF��������O/����O�]<�|�VL�f��V�������_�j���窞T���Abr�����{⌡C��+x�_�Z0C�?�(?�3hi0gY�@v��qJr")GDesJs�׫������p'��b��N`�Kl�Wqi�{�����yړ��N':����I���\��u*��MF:%WN���w}�ETȴyY��ۻ�:��!�5ė�B?���$N���7ٛ�d=���8G��b��N~W��Z3�������$Ss������$z+�Ȳ"@»H]�.[79>f��	�؋乢qyCt�i�a��g*Q�V�nmPb��O��3�D/��b��q�QlzU�_0l�˾w� �ϟ���;��G�&��EU�Q�U���S�FMm�R�5LK�c��d//W��*�䳞�|�6 �@v�h�|;�#�<<�ahz��X��i��ʡ��]���e���r(��\�)޳�
��đ�Q8���|�٭���1��yiH�� {��;4��l����`T.� a���XY��F�GJ��%�4x�܅����2��՚1��{)��X,3�p�nAjP��d�� Q^5|R~ޙ9i5x����<9|�����77*���5Op/o��S�y�C�R3�~���q�\� 0�`�uS��6�m��D���_n2�h�M�s b2r�t7�I������S�����g�����k�@4�Gc�uK&�ISr���ۓg��U�c���3�@A�q�^�� `B}c$ѧƈ�j���sz���Պ��Ԥ�Ð�b�?u���B���zXj$_�{���sڌ�`��iO����B�IW,8
)!�;P�Կ�Qku/D�&��Χ�t�E��C)8�5�l�|�оx�9*o�r���t��$��%v�b��pޱ��qy�Z�XT����+�+�!}ۺt��-h/�^y��jS����(1����[�%d#�����z�����9�W6(4L/:�p���+F�� ����˦�G���$l�<�IEr��P%�af�LE{�Vp�+� =����'���0� �.�30�$ɕ6P�m�mH8}��;�֨��I�c�Bj�EFpI�D�@{��:hg�-��Ff�K��Q
0��$Ƶ�^����&'�d=��t���D���?�������F:j-_��Ȉ�6E�
�wӏ]4�y$p�M����?��\9k���w�RLaL�,�RaE��`�4f\�Y��,�џ�w���ΊynA�7րC�+@4��9�I#�^�����/�]����RAhΛ��)��G�� V![�X>����穤�l��ݟ�_W�j��u�L�s@T�n�k�*��0��p�8wwx�k1P������\氣��A�	1pP&ޘ\	�?��6�:͐���4K.]�&���1��3��,�N���B0��g�1�������,���@fZ�#��!^~�5㹁5��;	3ޫ7�⬖O��w���">�L��Ii����J@ wk���$���C�H-�?emK��:��J~�=;��\�;���ቆ�@/�Ò#�	�y�n�^��K��h|+y�y�i��ٕu�lY�&�g#�`ۀAŠ�:m!��U�S�6�	Ca��;�}rg�Ҙ	G�k�_6��Шa�\/�T9(�I+kjC�J�M�&��xG
���F�"��?�J~��/0O�Q:�� S����	H_�^\�U���;AV�̵U�T�Uf���Iz��2����IC �v��lc]A��������O�Ly�C�P�m���T��2J�dȈ�]���������	��)������W� J{,�J�.�ʋ�0Z�uxB�6�4�mM �z�3��q/κ!���7�2uyj�⒘����`����ƊiE�:��U��潰SynrG̼�q 	/�U��?芘�SX�5S�w��Fp�7g�(KZ�$�$u,B���D�h:ۨ�'}CJ�H��_���UN��5H#���8>�]��y��d ��+�_�۔�k��F��ߡ�'��JT��2<���s?��o5�O���iI�j	
��/�s�-q�sN{�5�a\�l�&L�3��β�fb�q����o�􁤨�h�h�?� �0��,��p�"�{� UD��f���1��M��a�ܳ�F/
P�����/�=0j1����n�Z���JI��N�ם�h�0��0(?�]
���w��E���o�VIڋe��%�z�Kn �4i��]A��Fz�ΓǤ�-��+�i!����|\q�w���a�
!�89C-�piNfL�[����Tй\CK-��Gy�p5����j���������i���ka��7��AJෟS�Qh�͘�+'����M,��p?mA�J�W���i6����G�D?2H��+�G�&,�#5p���r�h�� %, �k>?� �k	a��=ba7}��C�!%�NTq����?��"���>p �>f��4�a
@��N?�A4�uB��Րc
�z�$�A��v�(�=;����p��j��muq���ԅ�"g�{4�����6� A5��#y����c+��x
t�F	%(�c  �g�)����P>�P>B[q	b����ٻ�ڢIZHHG�ਸM�}�{��\��;h��-��imr'ѵ�u'�����]���g,�\�{V�9k7�m��kMs���zYVѰ{:.��ҍ�pP�;_g� �u���=>;Ǆ�lHY+��O�L�PA1�oA�P�2FIgv��5@�I�T%s�8|���z�9@�C��+�o�KPF�UKO�38�q懇�8!���M��`��zw?#�݀0�4K� {.W#Y���ΪGi/�^�����Ώz��ZP�W�d�9+��`5��F�_?�����l0\c� Ɏ»�`xO/����� ��FU���䌩u·�ݎ�tH��!��-n��d>�X�dj��i���ەz����ה�LS����D�������][(ң4�rOF��Fʟ/��	木��0Pg�M����D�~���L��B%yH�*J��S`��ת�R8����k�G�:	Ĥ���:��i��ܗ�d+�z�W�3����N�W�+u��b��[��ػ75z��}�f���v����h	T�/�J���d]>p��+���.��1��鿐�v������jA�q#��]��Ͽ��+�^��Q��%�l�`�� m�-��hg�(IGo�&Y��=Y��>�q�a#�Xoŕ�aC�I�FgGٛ���|�̹�bT�ձw�f�������Tr�]}�ֺ�~޹bMe0)q�lwb[L�.���p������TJ�m2	�����2����Il�9𶕣Tɶ�OZ�~�	U1�����`)�D�A�Q���:q���q�bD&o�[�<�f��w���/�vw��bw� �O�����ny�9��Ł�4)yWèU����� �H|����zlL����ρ���Cb��=���5&`꼋oAS�����4�_�^gSXkrI'����!�7���o����r���'��a��됙���^\ +�l��#�f#ž�úbL��Eoh9��Ic,鍩Q#��z ܽ��l�҈��`��E�R�u �{j317��K){�'*}_�nq�wg(��XQ#�:�����t΁��+���d0��3k�2"��*	�����W���s/�M'3���>�u��	�J�Ҍ�[�Kt�HL��	"����_X=mo�@�9S�s��br4]�� �A�v���4<�� �V�A�����=[: �e7;S�y	A���뽗�R�['*�"xG�\��>i�k!�'��q+:%&��!K�i�y7N6|�h��d	�rh	D�5��y�"uRm!X�����B�IFj�n�CK�[���鷲,��uJ�Z�B���T/�����2�2��K[D Ț� J�L��p�ɻ�؍��-�~��[j��"�#��V�h��B`"�c�c��9kZ�<'J�}Ql�G��=a0�sN��)��2#��O5���6�u+�ì;����<�E�	>������9
h"L.q��%�ķ�
fpӪ���@ܛ�+�����{��u#-�Ѓ�8����U�VJ�ϳw T$![�A�,ͥ����7`+�y�農e�4-��TQcq"�u��ql8�ڞ@/����l,[Y�\)�1�;#G�%�"�[�J&}e��_[�ϱ�6��J���&_',�+v�K���$�ysJF.�m����i`������ʴV�Τ8+�GgI���J�M�>�l=g�)�y2���"2�2�����Ϊ�_F��m��#5�&����'�"�����I���J���u5�O��SF��l��ű���%õX��x�qN*~�"��	�Z��ILX[s"=k",�RkC�]�KS[���|��]:��)R�z3��K��2>��!K`��<���˹[�3���WrY� �����^0�31�r�t�ܜ�!��1��g+���m{� ��+}��E��>��l�
�7A��s7��wS�Ͼ��@`��4��ݘ[��8`m5������Y;��4�������-k���*����ړ�xs�ޅ���&�W큓�	~�t�i;m
����P
��i��@`�e)!A")t1suz����oz�r������K��mX�
3&"����q�����gD�\��L���&η5� ,ғ�e�
,�+bl�Շ�tw�KG�BATi /P��L~}1\�Cp���;���`2AA��%<_�d^�'R�h�)����Q���!���ؑ��S�R�����a��\m�7X�+
���|J�B�>wҴ7�����+\���$��q�9?q��"�xv勦4aQ<����[@�����GW=U���ǫ*�>U�ձm��?�?�2(��~�v��N�̡��Y!����>� �U�.�K����z;dH���m�k��	��K�œ8����(n,�j�&^�5����/7Zy���҈��>φ��fZ:�w�(~/�ข�8R�����v�5i_�Ŀ���m��@���%Ys������9[����F�.\6E��ن�,��<G����h`��r�z�%��
#�G�+�Xd�(t��/���a��CI�层=Y�$���;Db?v���:_�Y�+����Q��Y<	���qiGB}n��2>-\m:K�_��kN��e��09���ĺ?�mqz����mY�,��_$v��@���*��14N��R����AGOn�DT��T0B	�7cv������.K,R\�^p]���xr�6��w��E!��g���}��-f�e6���?��L^�Gil��uq�Y#b!�~��g/�$ �5��ɽG����J~��)�*��]�!�T%�38ջ��^�0�#=Nj؆L���۟a�9că�o�a�k/�y4�>Q��Pػ��7��������'#*VY7NAʙM��"������]Jx�oL�O�F�2k��q�� �bp¢�}0X���q�, �%�[r�+%�xY%���k��s�<P���g���ū�9�Dtj٤���bj9U�{�t�yY\IQƕ��HĔ#'�j�Ɯ���Q������P5�;<�,&1F�+Fܑ�rDƟ�bG�\^^I��q^���D�G��[���ֿw��D���U�r�F1��=@<�x�)Z�w�Gƍg��ۆL�"s�(ڃ�5� -���Gu�l��}����E[����L�J��nS2Ѵ�����Tb j���8��G�	G`9��4"�E��EK���$��n���yH���0������{�s��"��%.� u�@k���qI���������80�K��Ц\��} �j��	Kd�o{,���2{t�ye'd�u���l�����g�V�TK��T;螟!'1Ƈ�_j����WN�KHF�]��E	�<�ʴڌ��[ځ�<���X�f.o�YȽi�L��Co���hd��s9���5�k4ڵޱ�
�i&��|D\�)T��eR�����$��Q�����s�ŚѰ�+G��=%VJ_m�oUQr����s3�̻T�� ׸-�d����GI!�;��a�[�,��-�qr���~�`��*fϩ���$�P8d��u�ŵ4�M�Dw�y�e٠2��qn�ye�M��8�?�&ԭgh�b:��Ň�N�ʰ>�nK´�7N����!�<���ѥ�HgZ����u�'1��"���m| ��� ��x6��jܔ
Wԇ�ǧ�@Ƞ��$�Ji�����QFd��g᫤ߡ�vی�15�7��)�������#5!̶+�nD?��[�M�Z��Hƈ� 2��#�f�MO5��\r�E�c�ib�%�Ja�΁��Y��B�1e4x�Aʓ��o}X�/Gܝ���|��=��Q
�Xt�WWF�/�<K@}6�Շr�,�_mn�ާ���_���
܃v��t0���'�`N|A�١�����9]����)���w�S��~�p�t>1�9�w���JiZ�[�|�T��S ���I�eR�<�0X@Pң{_)񨰱�A�sp�8ҕf�S�,]��ab��Ɯ��׊a�|���J��[�_�&�:Z�+R�b�ZT�'�X$�h�N���S���bB��g�.��_���+��[ $G�=�׃�T9�Q�E)��?(�|��G����T�����'����Z՝n
 XDW0x�Y��ĚD���s	?O�>s��E��4�T͡t�]�����o�!��mEC^��ī{���%������ M9?�)[im��$�٣se��CT�ݏ���C?�Q�(���E�@WՏg�5U(�����d�Tb*�!)Ea��&v�47��g�|
���9 7�,]o`>.9���a}�i�k&2�qV�'�����vm�"n20��ih��T�B	U�Q�y�#�$؃S���S������:���Fj�Ev �T��X5Mܹ�z��G��ɸ#����$U�
FXl���+h�~� ��W��y]|�)�M7v�4�F�MУb�pb$I�5��7����j���~r1?8�Mb|(!� �^Cb7�ϟ�9�e"l�����?���f:i�7��փ�$�0����0ਸ$!�mR>MR$ջ��]��o:�X&O9��6�i�	?��A0R	Fe̆��£���=Gs/Q�']"��haI�-��vƶ��	7��b��� ��n��~�7������Ӯ�-$F��eh���∀[����8җ�I��hLO�=�yh�i�L.U��+�	�ϓ�H/��������]Beb��M?�A)���o�W��҃���+�s�^$�'{5]U�B�]�v �єqv\�@l��Y�M��
�;(�A��^t���uB[H���x! �R@�,�"���OJتЮwsF�kW7����;��
���L۵l�K�F;ie�Ne�\t�mb#�#/`o��k9m���*ΖX���[Λ�ec}�$H��.����Pkg���gT����&M��h�|��'�J)DQ!{2��io�9jY�xb��
/���T�I��ȱ��#Q�;*Mdv�_��+jF�|���V�XU�H�#�?#Y�O�=K����/1lnt"KwY
ۇe��y�Y_�h�J��ՁN	s�DlM�T�t{2���(d�7�k�]�dDS������4l�N=ܹ�)϶�|Zo�Ia�� ��&�u�ʕPϸ'�)�p˅N��}�gNJp��wͼC��+�K��|]߶-@����P5�c��y�<0��o?�kI�Ƥ�ʍv����1���MAE����^C��
�	c��_����T3��e[�I���7S����p��s���`�z�ڤ�O�8<X�\`�Ya��m$����N�,�Z��1��d�n��0�9������"�k{i����M�]o�F���~ÎQ\pՖ����ݤ����:�!sOtpB����nA=μ� ����eHfi��L�ݟ��`Q��He��s��o<S튬dd!���&!3LEos�mޭ�9��B���p�T!)�.m7��5:���Q�?� �P�~�ʮ�<��q��`8D�K���N������a�Ӛ�a�.���Xn{��z����=8�"����;a�0n��
	��������00�)?].}�E��s#S�X�;�z�ƹ_�z5S^�v�����d��+T��0=0��}�K���(�B撄�uF�@Z6���V��p@�X�'��b���,���|���5i�A����R	F�eUDd�݀ӑ6D3jV�����%���5P��!����)7��F"m̨�m8`���˃���Q���ϊ�JB������Ð1fb8�O-{Zi��iD�ϛnf��-����F�׼���wbP`z�.��c�F,R����"vż����A�zA��a�)^��L��<�Brk�	d�<5�>�\�^��n�!nrg~����${�v�p�g��}Z-�_֨�L���?����h���"�.̈́}�dhU���A���P[���0H<P~��l��F4W�|ӭ Cz�n Ị� �0�?�?1\��ŗ��U�I�7�o-��UM�t�vM�l4��6�]k^pm;	��y������PG���f����c�]֢��¾7֤�#�,p9{r�:�C z	"�>X�- �C	�ש�����*�~w��j#̺y��ͷ�itLS0���m>���Y�a-�ewBB�J�t��XJ��t�"��{������*���*P(���WZ��TW�">L�v9�'5�D�Cn�"jC�s�i�;���QS��^>���#ɓ)O6�f,r�Mw	ѣcF�g�(�~�����n�}D�}�GƆθ�p�����nFn�ǤL$��oj�Ѩ�,= 2�~>~G QlF��W��^�W�{]�����+` �qda�Ţ��γCQ�K����ì�,с���ڙ�eއ�'�:�.������0��,$*�(_����Y�� N�.s�W��Wɇ�8�5)�F ��p)h��Oe�[<!��wDy��wӠ6g|�崧k#-���?f<e~o�Bͬ7�m�@����P�;�M�~{�s��cޜ�S{厌
����l�G5�H����o�- >��D�5i�Y�v�(}|��H±�}�ٿ�H
�F��g]�?
w�(�>����O�&���#@.�|��#���kQ�����wa��unכ�>�$ ^��G��3yVù�~5�� kHO��6�{+�x֓g��&N�"q�F[a��׉��u�勐E&\#�ْ�J���A 3?s�c�x�]��b���l�Ʊ�}�,�.1 �eqF)BJ%Pֵ�<��z��j���s3�����<�iƇN�$%�>��`%�]��`�-Ћ����3C�k������h|V����οZ��x
,��ƅJ�S��0�����:o�?�&�v3D��f�����AO���X��@s���s���A����&��(o��1�w���T�t�ι:�A	A�5);��
W�*���9m皋ڢ_v�j�>L��OM��Q,Z�Ou���}�{��<��������F�� �f���I
�2_��|L��'�P8O&�;
PQ�=Of$8D���ͩ��-g͇͑�!��ie�P�
a%��:S�&�f?s�!�~����ZPg���k8}��V��K#oBF���G,�*}�����iV��d�Y���bk0��p��v�T.y����t;��e%!���o��=d�V���5|!m��{��}u<���y̜aV����H�V.�}((��UI�CbL��TG~���qы�U�WH\\הx��D�z��e*@YWsH���U��C�4P�g0�;�4��ˈ�w��a�S��ͫ���1�ۣ��i���+��F�����ۗ't�G�66��M@�c�g4�K@������o��Or���ʬR�|�r�y1��9�?2��:6�U������Gz�62г�g���+LX����s�7���N��R��v�ԧ�D�,"Hng
&е{��sV� j���<�ɕ 2ڹ`y����l-��R^$�<���$�r�I�9�gGH<?����5�,O,�����$NA""4wA�M�����	�Iy��d
^��� ��<F�`(��a���ږ1ߤ�2ϏQ�gq�ЧSw?�9̋t�^�{�E١��-q�]���Y��'�;�����Ń�'@2ǂw�CY9\Se���)��Y�o�4Z���=6���s8t��)�'�p	̄��;��Y�w�ϸA��C)�Q�}
���i�����幤��5u�"�����E��y*/㓭�*�y�?��TmTI4E讀� Yr��HG�?;��"m�VS����l�C���F�S�_���Z��ן��3���(KU&�>逄%�	�B#�0ı�A�t~+�����?��ćZS�up�*]�¾�#֌+�
�6�%>�_�S�}��K��w��V�����u��c @�uI����@^Dݽ'Z��D��V��;�+`\<�C��8���j�63��Z4%Ԯ=��Lh_}9� i����*L2����f��C��},7%����m��G�
�e��J�!�)����f9E9�5��`�-e0��u��c~�`F��C���&vf1C�B�s�:'l��ý��M����4J����G�>3ɛ5��G�����"4m58���l/1 �8����ry���������NA�>Ǵo�:��{Vi�pU�ӈS�Λ8��b��_Է���qJ��f���]o�x���� ^�i��c�e��0���S�lʑ�.0��Nv�KRx,w���(����NQ�dk���"W>TٛJuNA'"�2��i{���a�|O���A~�"t��ƇՀ&ݠ c�}��V�����&-��J%b��D��s~ڷ[�ѣ�P���,<_S ���c��M�nJ�`|���NX2���u��V�qK�F���P��/��|�#G��_�6蒦(0P&l;ū�3P~t� ��w�'�a˔d�s�9o)�6�Ćgq��T!���دe�*�汷S��sω���=��62�2��V�����'�[B�._+����ť��Y��\*q�R��{s����:+'������1���լڠ��C���G��&Q��W�(�1�3����u�W�G��مT�#G��AVm�n�a��*���q��3M`N����-�4���FeP��"H�hSqI�҈ڢ$��>C���D���0�ۨH�݉hU��R(���w�^�Ď����3W�Q�.>�R[����5g�0��3v���Q�ů��DB��9��C����Ƴ�Xx�(>D#��ܹ��<� ���+)�²ɴ�c���%:V4�@݅	���+?�,þ~0ݰY����뫮K��v~��!��iΐ��1%=�PQ,x=){�E����b� O��3�/(G�8��9�4LI���*�Hn
��l^/�����CǪ�C�4*� G�_�����h��ϝ�Ӣ��r8sI��WP@��Φ�}ɢB��	�-�tn�o۬���G��r�G��5s���9,������W���5�1K�6�Cn#�7_ ٥~�L�mMi���?��)��5�u
/�t�Z�*#�<ŭbC`%\�6Z�`�UK��Y	�T��sn3�-���8c�Myf7l��軝!�m��G���V{�����A9�r�/�fE����<XK�����R�#�E�(��8o�o�i��C%Ͽ�'+����V�,�
����Tgk���J8P����F�
����>e���f�4�F���\�F�5_�� `-3�C��C���!��:3��@�k��:�4�t��8���?�X�a�c��h<�l���80�<<}��bV�Z"�p~�A�)J�����::��?���W3 �����%����ȽG�sBW��'�f�o�.�, o�z�7�&B�.v�&@�����_�����J@�ߥ̲	U�e�GGCV�0Zv�P˻����-�Rz���T���}�̴��|�L����B�M�a�m������j��Z��:+��f�h�Lo�c�>k�?Μ?-��'����&-q<�A��1��u8��@�Mr�Bn��{�#�[��3X-#��`���rJ&�f?G8�-ĕ2|�Ř��U�|��yA|�O�j`+��̊vz��V�M�Ac`�f���7����v-�Ǽ�����r,�&��yǄ�-g�">RC�ƒr����lZB���(�q?+s��|h��䆲�����-p)ӎ���Öa�ݗ:�D����]�o�2�ĺZ;�����4����"����^�|��K�D+���gǪF���u6���}+r ��D)�S�y!�#�؇���X�%̞~�*>���y�e�B9�w���zV۴��/!<^��'6&��4��0r1�/�pPg���;(�:&�
	{S8�b��F���@qǠw����k��]����B�𢗙:2�����2��C*y$̋���^��+
zo�c��ނb�9}��z`�U�.m�7e �ev	���g�a庈�v�d�XfdGMx`��F �`��2����?�4�4G�¦�Bܒ��n�hj���ĚD߾]�G�8:0�Sr���*`H��?�M�ծ��D�i��C��Χ ����z�a�@��;�A����~Rȱ��Ccx��� ����"�$Z��ۧ���o(υ�I��S�~�!�������h �5�t�K
��-?q��bO�j*`
QbL"?it�9���,��vp��n̓�`6w��ߘ��UY��9�^�*`�l�QG�� � q���Ч͠��m̚���;	��ny$���hnp�O�V�(l��o�PX��|e����{z�e���P\T�*ꢕ�{�=����F�h������^�~^���>�m�A�5�AH�����m����s�r7���|Q�v��7��/��f���Ԩ;����J��<�GK�>˵��u��4%�a��quh5F
���\��*)M��O��d�X��^B�����Xg�Y��~����pv*7V�<\�6yH��]�s`je��e��w�N_.����#R���o�a���Hr��^����\��*�h�wV�>�d(u5
@N2�~]�AI
®����F:EIH]Or�N�-GZ\�ʊE5Aeo� ���,�ׁo9ǮbA�jL�,#x)� ���c��"ij��#6�5c:���S��eR(����B/��|���?�3B�t��#��N��T�@��bk=��K�/a���]-&0��U�J����
Yc����@κJ�(�5�E�'��x����v����(LP�9H>�O�DG|GE�%!u���24�qX(��y�gT�\�@8���a�ި�:�Ɔ�m����W�~�6fq�����U���#����mek�ٖqK�W���x}D�/(�Ã9+x�w�FŬ\���6N%#�#R��mx�%g����Ac~��+��N��l�艆��,��iu	� �.�=���<2�Ny>���;�V�Z���A��0J[�����qIw��Yě�k�T��l+��ݎӓ��V����a�^�nEYY�VF�jZ�����6�'�<8��A��&��������p�R�E���ρ�������ݗ��1|��	�"���R��%Qm+� s��� 
�5ON��V�n��빯���n{�N���ß�Kp.#���Dg�8���Olp�p]�p;�H2>/�"���S!�+���8J�1=���U}�`Je~!��ժ�*�񢖉v7�P�b�\0=�(ɟ^Xۄc}1V�B�
�����{��0��ު����O�[M'����S��z^~�|x��?�����%���;�C���ۄg!� 0��P&�709"����e��^�<?��o��L��PC7���@���:T@�d����%:�R�MT6��g?�M�����kn0�7�k�����N�A^m-�J��*��}#�N�Rz���|�U�Y��IJ��[�7�˘ީ��t�<�:ӱA�n��XRy��{�o�E�-1�JR�?B�}��!��`S˵��ƓT����%�5�jK�)�^$�.���OZn�o�8ߥ�#�S[��V����tO�78H�uϽ?�����h��sM��
�[_
����#�%:�����+�7@:�P�q�w���\����n�D�'���;�v�k��c�Gϟ}iiM��U!zƒU�{�Q�� \G�R�!h��T8�2'��!s�&�A���҄33m����)��߾�@fF����:���쇰f��,Hًu�Z(�a��r,FCc��ֺ7g�||@�Ƿb���3�PG��^��D��5�N�'�e`4LzS[����gZS��a��HD�j3k�5:�"e���Zr�׺���'�d���#ց:���qT�L��ǏU�#�־�/�� .����N�༻��>I��x����-Q�oCZ�q@���*��z�/��Ut��(����P�[҂�Gf��X&���J��~��u70=ǏUHx��8� ��Ĵ�*��(�m�����!w�F�%�I�-����2�A7�.�ݷN�GB��/k��� �P9�*_M��Kt�����������'�q�|���,����%�9,-lB��8s�Gϋc.�dS)�ɔ$���z���7� ���l��D��6��J�C�w:�����i�ʼ-}���č��a�8����U���K�8���?����Z�N��)y=���� ���"P7��9��lHm���
�N뚰 ���:n�=~?6x��1ރJE����jW��=�_���˚�Tw��ЙPIr��!5o����SK����R:�K���g?��FPk]�H�[��r�3�#�|���b�4��q��W+hs�]���T��L$�RD���ԅ�����&�In��xB�i3Ї�Sv����^3��p�O"J|���7y���������X{]�}�+�d��5��~Qy,>�Qw�+ڳ�V���n{ңW�=�1��T�-ףf��Ahi2��g>3j����+��l/lfe�������?�?^����, '��M���/Z���>$��`�|�J�JL��K�q�U��.��ۄh����t[���،�D���F�0J`}��=P;Ø��!�[��q&�2 �Z��d��r�c\��*���`��$0Jˡ��}b���&� �u6	���L��0�P\���v<v+(z�Cv�|��䨻� ��)h7�"p��˵q���%�.p���s���) `9f�rޗv�U_z}u���˖ħT��