��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��Oܓ;�������H��4*Z_hř@9R�S���R�:�̀T�j;P�AyT��[ŵ�(|/o��&�0�C�>ӳpo������uqcK�܆��ա6~��?��4T�M��p���Tx�1�:}wN�fɐ�a�~n{;��_�;��K{n?md�7�gi�����4<0�y���]aH�Q,D寱rJ�R��5`�A�{��
�;<K�w�?yN������G�(�Kw�&�uQ��6�g�'���)�,G}G
�IO��s��,��y�P��y4|�3�t�����A<��C�V�y�7j:���=��W�ì'Iu�}����׀f��=�����4{�Gu�eN���(E�i���j�N(�8~�ʏ�`�S��V��V2�ФC��p��؝�b5D�AB嬨��;�1vV"���?tQ��S�*(�	���im���}\�2�ijM��PO�y{�͜v]�{�2��\��P��*B��"��h�L�.����'�n�n�ٸ^9�8 H�b�h���K�p�!����B.u�l�V�*b&`ԚHh�є��ޮ�2ê?�m	s����@���D�ƾw\:��ծ,x�<U�SHj�ZJFJJ�[�WHg`�P����e��� �Ʃֿ�2?O;�F������?G"�%�Cq$,Kh����u=�$>�!�DD.��"o��Ქ���,�R�lb��wƬ�߃�C�8�&�W8^Ӹ;/�)nq2m<e���n@/\���L���x`�"C���FR{��������,�H꽣&CSrj.�A��F.0�{���,֬�	>gs�-
(1���
+�s]��$I�o}��6�m���I���`��f:=�:��i�7Q���*t.���W�W_S�I:υ��WƁ�E�"���|G��,��{���ڵ�1������	�t�O�\��0�KE��0�J�����|+al�|EcN����b�x����oӿ�|	/d]���-C�H(�Rg؍ЋNؠ��Oq^Pm�sJ1Z�'�����q�4ag��m�o:\�L���lS��I�Kw����sר�v��LW��Ƶt���R��~��+�[�{R�QwD�4!��E#�J�/T��4�`y�9-��@���%$:I���=y�s�WԄ��6-Hb<�� �p�3��M�i���V��Z�� ����%�E��N���}��I���a���ԩ#�;��v��6�ٳ|hAP����G�]�>�`]��2�!QM~��B��9�{�M�*�HV6�P++A�2T���)}�XveG��ו΃}��HG���_�&��i��A�Ps�8��h�\�>��C�m�	l�Cr�p�T���&1���=P�n��~���3`��;��|4�-6�豝r�`�0t1���k����rh�B�zW����۴hc"$<���e̱�h3$5�\����1���#�1�n���l��|ƥg
�U�5VF�kP����J�V�g�E�&�� f���e��?��Ӿ}���4��:c�j����/%2�W9$�14$��Is���xXMP����h��I4�#��Q�G�E;�%�٧W�Dn#4�
���PVjt�h(p������[C�i_� O��`Ƽ��c1�o�i����A������D�f���M��2�i����.p�}��]9m-��t�
�4���8z�����x�N�U���V*�b[��+����'�����ڋ���B�mv�q��U�h����b��J���Q���*� �K54bN&�����Gŧ6L\5���"�cm�}�}�	�3�,�*����Ys��^0��X&�a���J]��&qy[_�kȓ ����y/wעX���������t(�+�nlL������#�e��ж&���z��J�yVCߙ����[�d�#��<���O��3�	��^G�,���N%����ܗ8旃8�� +qe�����ƻ�S�'2rЫ� U�_��]��ǧΏ��Fxa�Q���J��ϓe��{Cw愗�M����r��?�.1�{?.0/
q��<�,z�m��xy�{�琂�Õ������|��N����+R�.��}�MS��{�2�?Z��ET,Rk{�t�0�=�my�80S�|ZG?Vevnu�mNЬauL �:!��qmsvD�(}�]2¸�3PLk�uDp����m�)�1NS�E�Jju�W�k��.f�!�#�9��:�*�x�+��<D�*1h��c|&gUU�b�Z&y��m���^B�R�t���t��t�5�X�L{�w��e�2��L���X���/����.Ǉ�#����T���v��Y�ȉ
�����b�@�q4�Υv.�i�v���[P�}�z�<��\�wM�A��:�=�^i'x��׃|�{Er2�^��(C���&��g��ܩM�</OyyOW���N��4&J*FE��n�q������gy�M��i�憎���uԴV��G�=�@D��<�D��a��V��9�#�ꁆ�&�y-�.�*��4�{��I�%��ke�<�1[� -w�@s�P����gg��^���KZ��M���Dc���6'�\�j8�xU8"�(�PdH�"��G�/�x�Â��Κð��s�ۭ�P�ej��[/�N����=;�k!AVg<zI�CT`�z��#�jS{C�!��o��`�uG/4Т��X��ꂦ�&f���F��f���q�r��#�j�*P3��z�ꞛq�"�#v���4�',8�0B	+"�2.)���Wd��!�
&����������qN��j��;��}Wp��$vA�%���*>)�"�@��nmCul_���I������
�����aI�1��Sn/����8~��P���Mw\m[��"�v�@�V+��]ʚ�V�f ���z��oJAfq��lG����"�C{�3��n���o�㡙�1����L����/�H:kCx_�/ER�v9�㺖�lzg (����q���e�_�6tQ *A�W�PY�<l����+�����R'n�NWH��0Lc���C�W��r�Q�=����Wӆ���,Z�R�D��I`�Co�]*8I�W07pM�Z�O7|�~�-y�c@D ��g����F�B��U]GH�@�o~���>���D�V=�l�X�.n]��zm녩�1Ĳ1��Z�IwԵoT|�t9�-�h��TX	�*�Q�nZ�[���9��r;�m ��'.�[������j��AV�}c8.L�Dz���n�6hH3I�8#�y�W��@,"G��/X��7����t-������УL�S!���
`�]������XZ@L�]��>��s0A"��عo�OQ��������/&�R��k9Ό�0��&���'��<��Q_�\��"���YF
;z�GVN�����ӗ�z������)��-�b��](����8��@Q�*S��E�*y��M/jБ����c> 0ج�v�G,���G����%B��z&�Q6��ѡ	�@��Q�a��7�	,����ʆ����"����O�M|:�Hj��,���w͢Dl�*�٨B�P"�u���T�����ZH�-�����Z��6<Sl1�-)�(T,���.�3p��qyJl��y��u�nS�V�V�2�����+��b�-�ad�X�y�>$&���%I{���ͥA�M�5r�m�,0�غ"*n�ճzK)��e���_cCk�d�[VF�1��8,��H�e
��p^<���:Ze��O*0��DʂjGW+ȢS��ʐA(�����e�5�.��;&&�I�x��J�3@Y�A&�g�q���B��ʏ�H��k�`��
��ט�ZX���i���#����,%͗R-���t�畺�n���ң�@0$K��ۨv�ܖ�0�&�g�TT�������BO?v�-�ܧ��j�ϻmy(��0vd���@9V�1DM�
�5�H�9`���;�d<�?Qg�/_f��	�0��G�/qf9�>�3��&�;G�ȬZ��&.kΌY�e�,�9u8����NιDj��I���O��~+m`�O�!�����.�p���$�k\�՘ס�߹w�����l��4�8*�sʋm飘t%��%�& �{�zE2 ������׫�DKO��{�aؚ{@�>�m0nW����|��'������-B�RL+�=F�x&U)X��+p>�OC ��d
IL�R�����FN2t���Ʈ]��ո����R
�ֱ�������� �c`k������a��}� ���o�FI5'��@�<o�StCBJ�S '��U^,@��� - �#�+̓���/��������\�\Lv��dgu�����.=3aI��y��D>��ioqu�z�F��Iʾm�H?\W?y�O���sKDiCyN�>gDU9G�S9Z������r��Z�m����s�����J9�'Λ�(�o�{�nuGY'^��h2���qɜD�]�!��xd���%��� 7��|���.� !�P�Fe<����p����XI��qnJ�7�?W��R��!8c|�����`Os�M�ߋT��\� h�EX���ӱ}I �,Hqs���;J	���p��*!�w���1�K @~Nf��t��԰��5Ƀ��8��M�<o�Fkj>v�D�Z(�"����~��`[�-�18��{b]����g<,�� ��*j�1>�|��:�O{َ�1�m;�JFR?�<;�������4�QH��I���P��Z�f�jx0
����N�M0�,`��FB��3�na��t��Þ���	^yGs*	/�"��[�ȃ��K���y!���С���*�^���A���B�IXٟ�6�YW�3ܢ'�/��֦�s���s�O�5���RGXd�rXJ����u���m���m�#�!�H���d��zn�v��2�q�Ͱ͘���n��2K����?B���(��d��?�bC�̒��<�9��[ �`hձ���l����P	�x�{қ>��0��(#ɹ��킀'�8��;���D���ֲ���5ʛ�c�8�z���i��5��i��?	f|-�ȭ�/�A�ƀ�w�1��}
}w�\^�;���ec43V]#�u�:���:�����n�ـX��L��I�ǖ����27�b��HZ�9+P�7�uI`#�	�7�a�'�p�[��d&���쯭��������Nb��wk�!5@�{�W�c� �i+���w̱I���s!��3�#���=������_�B
ΝǨ���]�_��꾓��H�\��82G��f���b6�8z�.�J�Aǂ�vs/p�v�-#����
�Eɴ�O�1�{su�i�ԝ��!g����o�x�d�g=� s&rCV/����}_��.L�Ŭ4tZU��>S��	��y�`�-(�L��{��M7�>*�yU��m�$�� _p����~�$@r�yz����N�#��l�L�x��ͅ���5��ΞS恸����+�z'q��\}�����p�¼6�U�9eL���YU���l�Ny[��7L��'��VdDCro�v1�`��߽���MY�k�Ke�\��>��w.SҖ���&������G�"7���5ΒC�$�N�=��\%����kF���tA���Ѯ��6s�,O�ͼ:mKEkn��u�RB)���c�b��ۘ��x���D��t��zq�u�m�Oz����h[4"�U�����{F�NKk����Ք�vX�c��8�Fl������Y��^bi�8Z:���v�C��V�kg�pr��[N�Y���w�(uǚ#[�� �p��	,�+��5r��T��94ӫ	���M�g^we�6ȅ�
��Ʋ��R˲C�|�� ������D�}���X�Y����W�B��%@G�.���+;I`��<[�}��H��_�ޥ`2�u�{

��Ea,5�����m\�t3��D�����vu�����,�)=b�[0{b"t�Dl��.ٮ�e���1�'>5E0f