��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)�2������2p|�t����)D:�_*Z9C��]x�7 �E���X0��V�Q�`,PXӂ-�����鋉�7���U?Ϩ��h�\a@68�+#r~�o�:�Bi�Yr-x�d��@��`n<wW0�W���eF1"�9V�SA�>�W��L!�S;?���#-b��D��ө1��un#�;5 s����T�\�s2���t��7�>��-[���:�e�-��C��	̊.Y*�!92��&~�Yً��CJ�:�o�\�Q��Z��3Lͧz�ne�6S�t�p���Y��i˩2%8"��yW\d�0k�5<8���� :�T۸gr�wq�9���ݝ���D%���%�����W���K�~3�5�k���N��A��_Y��>
*�c!�^2��o�y�Bo��wzg�xk���]+���ȧl��{��G���bf�Y��v/ՌB�:�/����H�`��^���+bC����>m�2~����VI����A2��~ɂU��.��?g��,���o����V���S;��W�����?	�.��G� "�`�ܯuX��J��e[Sa����y�+��W2(g��U4�՜���S�mb�k,�\�P�X�/�	�>�
�E�H�W��.`Ά�`�#�6��R^�A�Ԩ)��x����x��S��d;�:�2�X=����"GI(��*[7�aA{J1���#|�F,�3�p�\�xyK;˔�"CO��w�B�ф�C�Tw$A�d��D�N%tK���
����)[T����\��ɂ����ʲS� Ŷ����H�(t<�?�ނez��X��9f��>���A	���ځ�/�� �Ć�niíX�����{'��\��r�W�Nu@7����c)D��򃚞�a��=;�׹����ˠ劁N�]�Ƽѳ���z�^�|�)�_��C��+e�rYY��)�Q@�7-N�@��L�����]�����֗sK%�t�M`�x��Եz񃐼A�3��4����8��U,n_��Y�t,���t�֑�O�)T�at"�B ��tt���i&���T������%[	�m��5�-��߄˜�V�&d����dXҘXɀ��d��;�����tnD[�G���n|�LK�|�n�<�H��֣,#�[Y�e6��"O����k�#���4n$�
s(�Ꙅ����Q�k��n3���e��O�"}�;i�m1����}n�=.�ϕ��Q������Z�	,?t�i9U�$���������#�i��M�X\٫jJ��rrU��ya���c�Z�ƙQ�+&��k|�����dR��&Ì6ںF ]3�d�P�)�"��Y�|�4�>ܝ>~��w�[ӓ8[>�Ԙ�p�ε�ߊ�MyG�B����䈝��?��b�ܝ�aQHj^���3��E�CB;U�0�J��'���_�`�p��M�(��轃��	#5�:{%[	C���z�js�z{��@9�ŗc�>��ᨏD��1$�����.^q��H�З\z,T�����J���:��gm�����6z�6���/��B� �L;�����P����ߊ� ��K�F���Ǝl8��LF��f��A��R�^�P~�����mv9����2�<�-��T���+�J���f�%���{R�.�B�`��,E ��q_y>"�''No�l:l�x��7"`�΁Ka(�(mʙ��	�&�u���	#u��K�����5G{����`^4w�G���G����v�����8RH�V���C�P���n�^;�6Q ��E'�T�#;��Q�L��8B�4��G�?�@���@��'B�, O�ؤQ����n�$���ɤI2i�J ��5v��㊆[�V^)�.�:��=��0����BҦ��
j����юO�J�Ɨ�5�5;��*�U'�t�"�"]�j�ž�OA�Mr+s'�O����+2-���/n����U�Z�Z��d+Z���3i����1<�O��pI�3�ŴS(���MP%��b�1t	��`)Y����id��i�P��,z'�2�z:��d����2�f�����$�b��_�(he���k$l��]G��Tٯ�_�rQ�>�O?8�a�쉔"�fo���J  ��X |hR� �ӬF��Q�:���ݐ�y�� ������l����w+�=J�>$d����+ĥcQ�ʴoq5�.Ž��b%W���׆��PX-k��l(�S����p���뚇�#'��%
,=��N-�@����kY�Vm�H}Wd�m�*j��T�����p��qp�]��Y�~oB��H�\&�	�|{�,�7a!������>�.ƺ�R|���)#u_���;cE���z>�f�j�l�Fx�a�Ƅ(y�\S�7=R\b���=�����|-��|����Wg�E�>��c���{����Ы@��1�K���.:*m��jيy��<y�\��ޒ& ��K� ؇2w Wԣ��΂2�S������t{Z��"�^w�uh���:5z��bc��CY�+į��(mIN�C��2_e�Hr��Q�zn�i��l_@���'E�)T���l�%���-W���0D�wO�J���F�:B.隬��ne�]dI���v�lz��Q`�4$h��b���e�I�U(��ǹ�[��5BFγ�E{ <�h���c5B��w��p��I��E;�2Ϭ�+ɺTh�ފ���%@#� -�/���+9����B�+���zr��ۅyW��Z2$��'�0[��/�{[�IR��j�sۺEDx�VR��i�V�.O$�#���R����N����7��CJ��3kb��=�\7)X25p5h]ͫ?��4[ƻ���AR^_�h!�"S$�[Q�G��X���}�~ګ����%3�L��kg�ގ���O�%��]�W�z9�/�֐�c�e����k���5�2�����,�agIpu�G��N�~��Z���^��`�J�6캻���:tY*<�y"����$�ũ��/�y�>��*�t�H=DP�Ά��˾Q��_���R~��+z��J��#��{��\#��7彏���Cf���u�B�q<uz�YB���O%� $~)��~�"��k{~���t���nxt��*F{|o� hs� �U��y�s��E���R�O����=~���w���"*P»��4/N��>}r�����4S��=�ze/!�O��:��G	���g��	�w)bz���!T$0��|f�\�	t�UY3t�V䊒|�j���ܢ4Ж�_W�V����&���^����Ӷi���L�2�2���f�J����֦X:0x�r�t��X�p8����w2���v�F$Sl���1O��4�X�)�i��|@og�}�ے�����c�5 �QE�xo�����U3�������K&N"�] Lxy�cie�39����K�r�ٞ�CV���r}��0�a����L?�	QgW��t��h�G ]�w�Xk�D�uu>���_��k]w��'����B�-�7:�Z?�T��l.
��`�=����v�y�B���<����[��Ԁ1H �Xg�����"n�撛�3<Eh��/����3�S�!�7YM����$�+i�7���! }�,�m&k-�(�v���iP��O8!<�C-77�v慿�ÐW���dD9�4�m�����R�x�t�{i>�u��u����������������i9� ���ؾgP�
����y����yQ ���	[g���O�EDo��T��c��6&U��#
�MtT��>����keS_a2�b���#h���z�ƺ��@l�>���c[�oY����H@5�K�Y��6�G��/iF|�u��&'�H�����j���s�$��d<�c@��2�	C�u��Jc0��2�|ْ.APf��S��b���gH�T	4���2���R[�fe�H�FƆ�m*Nq��ZPj��4�x=���W_�C�5H�����d�r:u�q.f~�Ѻ���9�;L�e_�7���4��F4��p�y��M-�s
5\g��o?���F�|�釧�<P���0x�K������iu1��g���ba
���9�*�^��=�u��3��w��*�?!���
U�>�¾�7�0��))��:��r��z����3�{O�o�Xd^h;�s;�BO����t#R� �<Sf�f/�rp�m*I
Ϸ����W�H]6�=%(Ws�V���o�a���ò����5쩓$��)����ďg�,������G��\�@�M�dw���԰^�h����?���ׁ%�;8�2��fo��\��HqeJ5 ���L�9�D�Gp�w�V������}-!��o�4����e+��֘sB:w��*M;Q��fz��&�<�Or�ؙ�.ғJJ*�����t;��QBz�/nᖢ�m��7��xTd��qJ?�#��`w����i:ցPԬO�������e�*��@�����Y����뜚�70�7��y�������e�ݪ������]8�T^�u���Pn�u0+P�>�Yo�0h(����{�#�U�jt�UkB�$jv?SuW��2���D�-�$sm:G�HJ� F���O�(nyO����=ĦE�S�&P��VN��ͧ��)?��y]�CZl$����$���+Uc���IJ �M6+���4*�S��%o_���{4}#���:K'+��z@�)3�b��:�����|���2B�8���W<w� 
y�jiq.�Z��������h��ݎ�.��2�S�Bܗ�����g�l�7����q�i�7�|�k�����W6{N���U�c���?�&�U�a�>��J�
'��ZSu�f%���(�ٵ}*��)?�+k���g���#B�.���`TKeWn���&%�%2�X�/�����oU
�;���f�+�lX�y� Q��zC�}�hc�5w�rp��Ř�{Y����K.��j��]g1C,����v�� �����eHl���,���"Q��_C�VYg����c_,���\�~/E9׻�=�V֋����t�����Y������_`�E��N���/�xS��)7�=�����.ܞh3�ANԸ��r�n�\lzR�W��Ȃ����¾�cԬ,���o`� ���!�sdW��b������$���(w��_�ը�+�|�N�_���'}3�6���y2�5E��a5m#;��j��U��$ѷ�t���_�j�F��k|��){����}_q��^���3���	�����?�)��e� ���q�[��U�8��N�S,�Ѷ�q}�n<3BW��#� +��~b���r�QV�	�4ED�QF�m��j�'�"�}N����`��Q�?���v�xl����Y�������3)���ez�券�JK��/^`�[��ˢHM��ɕ 0��M�-p�v���k���G-���"�oh�Y���:�'�m�������ˑv�/����2/�7���8�&���+Y���/K���zP<�t�����C��N�����B�br�ؗ���i@�Rjz��9H��j��,�|F{�)�}C����J�>q6O,�.��/���O�R�_�p����� ׆?<�bo�E7�%_A�O_��� y8�f��e�������uc�H�1\*Y>WTD�(PtE������j�G?���g�3^���M����(t��(��H��Z2�K���V'��@V4��3i�X��D�r�c��3QM����ve�?���1LVu��?b ����K���}�����y�_�k?�/]��ә��si9�,�xjEzL��#Q��"�'D�J:U5�L���h�Q�R ��6k������n)6Ҧ�N�F��y9
S�25�̆A50�����2ҭ�S@h��2bK�K�����=��?z-�XiR�lʄ~a����-w�!#��"��7x�ߗ� ��b^��_H�mh����.n����T
���O�d(Qe�DE@J�&�	�B��*��\��P=+����x���,�9b���t]AH�ss�a<*z�3�C~濥h��TжYp_v`��s?�t!.�"��٥π�<}1'3�Z2X0?�O� h��Ո'�����(!.yE�TOx-�c~�0Fޔ���#�/p'=�yk�tٛ5�۵�������2?��gz����T6������e�}�-oP��C3���bep����|�5�e�~��3]9��=����^�!P�y��n����ƒ 5��#c��^�/7ߛR��,�W���-��h���tBW����|>OĈ���Rl��p�`�Ah�N�2�e�Rl�/�P:������x�A����U� ��ԗ�k��N���2�*��Lܸ��w�*ߒ�9��h�	H]�7��u0V�,2¬L]GOf��'��lU.�͜�ұ(4X��۵�P�*��=�m�q�@\�˿�U�m��҆@��-g�H�M�v�wq|�`��=�ӻ��-�ȁ��"%��:��4�EN��ź�T��4
��7�P���I�>�}x]��\��Y�i{6^������n�ZcG�`-�����1k5���E#�wl��A�iI8�&�^��)��-wP�)�*=ǰL�O���Qٷh|����*eJ�D�6��D3�waˣ���h��W6E�^�7�G�6;x��tS;���m�T�.�;�A��ߕG��w׼?�]4���b���R���;�'��j��Z�8=>�@Q�,���{����yd���&��祓�U۔��|�Dv��m��:���� ���#����i��_{�]��wF&��Oupb�S�\J�G�)�+��4�������/c�-��V!\J�t�BF��
E��]��K0��-~���!�v-��p[�	1;�o�q�"�֚����|F���\�*3Z��qO��DB��q�	�'��:�f%��3긷��1��bU��j4�֌���؝�F) �d��Rc`Hm-�T�(�����S���Ob{F�����r�$�~���Mo�~�v/n�z���Ok�PP^˜%�z�c����X/��,�rb�SLk���7޴��"`���D��bqT4�����t��ؕ�z�����Ѭ
+�����JKi)?{uSb�F�ז+�Þ�4��N�>�.��:��f��؂�3ibF�P���q;����m��(�~g��82Y�����. L?�s��
fl+͐U�ԓ��z`��2�����ع�au-������Ćw��\��!��=x��L���j�We�i3-�A��LD���(�i<W�ɸy2�@L��7���[�t]�=,Eo��ptՂ� ���?����d�:���g�͊0�sri!�e�(HJ#��Y�3��}O5�ʵ�<�a���y�FtR������g��}�M��s1��;��o��N2C�=H�P/�_���+����� �d���(:��q2q�A���_�w�`W$:��Ep���ߥ�Ƕ5+ z�h�
>�+�7y7S%��'�"�_��o�P�+A�:j������=�z��Z��H����/3�Z��`Z؃zG���k��e�>&7�ջ����K���"trF��,�M����ץ����v�&d��1k|WP��ZW,���5-�$��0�9���9�Ld��A�����%|
�Y�?�~}���`�2zA�X��Pq�`d2�ي�'>�m�Q������$��a.�½$SCMxbb����Y)��O�(#X��N+Y�^�i`6˳0A7wj�)j�5�O���"�	b��o���Q��mu�0�gA9�5�s�4�Jf�پ��<ڤp��+F\d˟]�t��&`Q��z眜u���$wN���'~�]����Ї��72{ ~x_���:��?\�)�m|k6�q����=�O-�x��?����OG�oa������H����No5�ؔ�`�&*e�o�֑y�-��De����.��|Z�{��2���6��8UKoF�|O���������cMl���˶%�?�m�Q�=��K�D�@%�o(��`���^��	I�#������'�;�����d��|�􏦆�QY���z��&
�U�N�}E"�D;�L5c�p1��[\���%�7��`���֍	��Q�u��ϲ�w�����(�5pV 0��q��	���٥~a��"�V�ǫ���܈��A�_�;TQb�(��Z��T��zI͋l�B�w��[ے��*�F>vꍇ�T�u��'F��T�˅5�-1Mz����c�W�)�����`k~����:��A\~��MZ"h��n�_	c+9F@YVJ	�t�M�R��oU��B�J�O�q�ڵ����� �.��M�Z��z�Q#V|�qj�}��ofP�s���^�W
���=�<�n�V!K���J��u��ƊD���x�@��$�5�=��FI��Ֆ闕*OSV��N��~!f���;͕�
9�A���̀܉oƣ-���u4Jȑ�A��*Qj75HW+�T9%�i-t}��p����2c�=;�Y-p����*�`�h����;r��$�.1�~����1�t��ɟl�=���T��F񅧥�\��Ə0i�o���	m��p�w���&���x�����s|]|������ � �aoL�N���}�������kU�Ԕ�"Z��q���$�Ղ�N���-���<׬?�t�.M��2��K��p�dY� k*_���u�=h;DYJOҍ��S����hh�Zs-�T*B���NQ��nr�ò��E�U\�v���&�_.Z�Z�4�|���$*���i��?GX/"+@�Qn}�F��A�c3c7�4�P��?H
Z���1d6-�+���kE��M!�{�f��N���;{䄻V��}�gQ%�͚J��i������=6vx�*ĕ�=��!��+���[b/u�����e{�\/8X�(5K�A{L��H��]3X��/̈́�!R�2�c�$>��?��Y.��Ȅ����b�;�B#��5�cJ�,�.���	^�.#��+���m�a�lz\phFP��� ��54��i1t:Ԟ�O�������P��Rv�A����p�����FVz�GQژ9�>��k[D��ݛ��6@�E����s�����M��t�����YPx�=�����$&�����̹j�s�8��EF�pQ��\�^P�阕>2d�i�M�*�J蒧YŢ�l��'�U��_���ā��]��"g椑gٕ�eq�k|��j%{?R��"�b���V8s�>e��PWp
��b� �ퟦ�Ξ�.�b k����;(
������G��ulQ��s�u8��&�6&�\��1�A`�1�=)ͺ�^�}�ļ}�.��G��F[�{Nr.�-@&0|�!x~[��}e�ǟK�����L������}݆��Xj�G�&u�r��ʘ�4�Q�]͞�ہ���O��q��!e:F�[���"���Y 
���5�<&�<����lѶ}�?���U�b��?4����ۛ�{3M�ju%�%27�H;Ⱥ�囨���	�/w�{!m�I�?'˱4~��tF�w�q���ϖp�0�S!ޯ�[��	�"��R����#$�eǕ �f�����|�E�%{�?�6�3�1�*&��I����櫐��J�e��?���N�D	"y�eЃqC>=�z�?G*���7���4�W��h�'���&��]��Ĺ�VVvHg^���X��evT`����h��=�ԍ.:�/�<w"�����k��\d�jN�d=���z�<�M�0ܤ� F�ݖ�"�<*VL6"�v�y��wN�՘��<f��jS��z�v�f>҄4$�r����/"�|;?����z�5	ָa�[UF�wAo���GԌk��C��9� #���������DIMI��y��J�)}
.�RA{���Ў~���V��:���鉂lH���40�VC	��M�F�^g'��y�o�X���Q�؋�-���b��be^�7�Vs����X8
3`��~/r@Wl�	�O��+�bnLZ�IP��J�m4SDq0�Լ|���9���#���p�7��ng[�v������B�'�O����ߋs ��ar��\9�j�w|�摯���n�2Èҿ+_���ڮ�ӎ�o��q*wQG�%{f�W"�Ҵ'8$�J��(�{���5?��Z4>봫�^���O��Y�0&�aS��i�E������^�Q�#�
��&�(r�xZ��S��������_W�^������$��M�b�P�X�y�MGfw/��"8�{lW����,=l�T�F_!�[hU�]Q���ү�gc�p�q���M�$��y��s�L��c�� ڻʜn�0������V�/�t���V��A��k�b^!������M���ed7:1}�����	v<�CS�oőX9?����e���+n����Ձ�v͋o B�ۈ�oB��"BC�Zs�q�eyC���+A�{(�������(Q/$ͥe�r̚���ܣC��vO�S��`KN��FN7�>)_?������a^���.)�GX3V�E�A^Z�f�">N����~��IdRR�苁��S���I,�7D�".����D/8e����)k�O6��P��k^�җVV[^"(M�ٕ0~4�axI�B��1�d�ˋs ~딠QE^�}Xn�p+g��^�q��nҙ��׻堭���J1񶋙`Z�d���p躵��������%g].�Zi�6F�q*��!i쎜:Y����FI��#-�L�G��n��#���Jc��S�n}l��D<x2C3k�Z3����o)�f�F�!{��I��#�M �]�|���#����^[c�{�㺉P�]oO� �� �y�T�&��bkA�����зqV���Ľ?�&��ů�R4	A�r�G�T.��K�EA�;.X�BB.Ҷb�(���ci�mGc's�E�%F���n�@��LԀ
>:-�����W'�;@�,�n�ٙ)�B%X�V �#f��D^�����!���T�����=��*u�\�˫-r�8�҇z��v\
�9(-�$˽FhP�x�«�
S."|�a��"�zQ٨����]�y�ȩ�o���ا����|m���K("%ӏؿ�&����'�a�w�{_��đV��^�f�J����@�qǴJ�K�оXڰ*xO1&3�ҡ�t�r7�A�Ɩ"N�Ϣ'��<wi:3�k������&��	�xo�1LǞFDb� �15�B��}l���Ax.
ӣ�%_ ���Fv�o��m�`�
I�,�q��{%�Ϲp�D`n;��2,�Y�<��*A��>ZFX�e��; ���eeR�lh��M>����mm����SafЮ3'|�Ib�\���t}v�wÄe�+M! E�y&Wx��{|9p��M�Β`5�� %����ԴĿ�e�o���}RR��.T�g��B��'#cl�DG/M��ӿ��JLD��1���VH4�������2�=� 3�t�������"m-��aj�xT]�e��ͱ̏|�Tz��Y<ı��5��;��Þ�HFzǈ��S�1U�i���a��7�נW���.��(�"�X4=fy^e/�r\��1�@}�[P��2�Z�BY_*h���7	jX�kJ�2�y@��
�_X@��	�{2a�_�O�f��n��x�44V��o����3v7]��+"E��b�K!�!��W�*���'%���,�hMd��Bn�����&C�t��!���D\��15���W*�ư]T��UK�gŘ�<p`,"�|A�ffr�7��7�Y,1s���������:�vb[hGRQ�� ����x���h$^-��`�,�3��R7=iEX���Q�O.�m���������#YƮ{i�U�OK*����i`�g�V@D�;K��{�!}qXk�l��I��	��3i^� �gSJOtF]���LZw�c�i�����נ2�+��3%��k��nCה�b��I�����;um_�O�ϝ����l�(zL´�"����ԯ�&�d�~fW|Q���_H Po���8����[�F���R�]�aE1A����"AC��I�;�����e���R��1�~�{`��^:nd�GLnD�r(���ӎ�qa�;�b3pŪ�q�HSe,�YA�D���I�7��:����x�`FcW���E�IF��O̽Њ'��PR{�i��E+��Ћ�~�ߡw���H]�c��t�#����g�ݽ���ж�� ��	E�\���ˌ�4��X��8���i���G�.���2�Z�8�G����I`r�� �z/E��[��Yu�p��)��=yjjf!w��~�b0KO��d�E�PP��l;Ӎ�)L�������'��������s��'�rE��u�p_
R���N��V/}�j �xE�RE�E���\��l���(�P/Ģ�wê]����W�� �)H��	��wF�^���8�Fj��f ��Ѓe�ԅ���G��F�X`�~
���GŐ�tz8���a" R��Y>l��"@g��+^��q�~K��绔����ay�F�\���Sx;�Α\ė������Y�F���b��ļ�	�S$B��x�[d�CWE4�'ڶi�SU��˹�.K�h1�*{�S��9zt�!M���$�0�� ����0�j�ǅO&�+�9W��$R��a]{��4џAl�Z�|�^��ґ�a~S�ŘSA��8
�쁒��ۚ˕ l��K
��V4q�"O�i:���W�U=�=� �E�]��w/z��DM�nԃ��g�v�t�l�U(l/b���ȕ88�D�w�3�b�� (:#�^���TN��*%+%	�q��~�@���.�C�$L�B|���)؜��*�8�ד��^�{wΏ�ER Ii��x�����)��*Kp#�FR���F��5�X�y1>���}q���Q�MTJ	�/����`�5Z;��)c�)��hڽ{m����(tۗ���k�p�b�vځ���L]/�r4y�-D/���<�9p)�F��f]y��w�R���	a,�0m��j-T�k�Yv��~Um`D��W��G��MP�#�q�baZ�^�G���A�q9G}p����>�;$��!��}���4.��m.�yg�L*x�v��
?K�:�~��e-��<ĭE��8x3����1>!jIRKԹ�2��]|�����`��@5�p-=8���w��8#E�N(�Aisd|cb�3<�_>�Wv*�i���:R�~���J|�'5���ח'����1l�J��`�;�4�xN�+��u^(���R]���g����e'dvl����b�A+V�`� _<�{�Ly>X��+�a�ӓ�@W�e���	d�b�}�h�m�c8ф�->��0C�D���c`A�-S�D	���"�����b�"�]Op�Epg�x���yIbP���.:�����W+7�SC�;r��=��!x�n~�%��&����#f�x|%�z)��5���lU�9.w�{f��ƻw��@�u�~�k��;��\���|���Hą�Lz8J\c��{͍�:GӮ��r6������M��x`"�O�u��jᗧ���;-���V��8�Cܶ���A�?(��BI%�v
�72D ���Ց+�)9ϙ,�F�1O�y�����^�QH���M�n�]btE����z�m�O����/y��n�Je�=��g��(�U��������;=gk�!~��+������o�9p�nJ��|m��܂fX@5h����`Ն���CGNt���bVd�C>�|�=�'�#:�j:!OA%v��S*�׵s�^U$5��T�����,L��2+�f���8����n�2�s��]�S���z�3���fM���y���`M����j�n"�W*���ySD&-k)�o����/��K8�31��|�i�_��I�
��;`bt���q�2�b}2�� ���M��`RI�������~��鴮�n$'+�j� �lw��i��V�գ�C���O�<W�GJ�e�~2�R��ډ�Lȗ�]�'Τ.�����e[�M��u�֣{�g�",Ӣ	n�3c?����̞��B��������HFOZ�ɽ�:
����5� 5���L�xA`�v~v����f�@��夸�
�>��ʗ�̩�{n�
��	}�5Կ{�n�t���`�
�G ��~P(�r"g�.ժ[�Ǆ�����=�'�6G��:�M`�� !�Tº�nt�a���14��y��2J�Ͻ����䤇MHq�hň<����bɠ�l�tG y�D��	���W����t��)
�w�7�R{Zk�qOʇnB$��"��22к�~�}G���p�+>i��i�x	��ej�����zHε�P�8G�c���b?�{���{��-K�LUq�|�
�=n~t9���}���%�=
{�&b�2�v���\��.�-o��(F?�����1�fa�ƫl��1���~q�쓳	(�w��n�%��x�����[׫�WU䦓,==[���%���F3��l++D!ʹe�GcΛ�^�V\5H�vwYv�4�E{!�c�oՂ+(��	M������BO[�͝!�(v��j���ͬ�d����U�V�7�u?�#�՝�OK;���Y����:D[� t��y��m��r�I�Ǯy�w�R�x��z�EW�h��̔�c@H��J 2ٷ�?�
]��Ӂ�F��2��:4!�[R4T���4^����ڈ�Q��*ц$�Ԑ���&�e.opOs�i~�|_��v[E����
�1�)1�7?�W�P�S�$�
�����66�l� @�;�R P"e���6�zw��ad~�Ǝ5��m��O� ��L�B�$��0�#����6-���ND?k��j���b��uU��Д��|eu�s� �����ٲ���z�u�V��ll�ɐ}1ߚI����$$l#H��̊���ݗ���,Z��m��������CY�Q�.KY�9��`�;?��Q����2Ŕ�/mv�u8϶2o��RS�������(��A�O=�c���;�Jh��N���8#�lM������d3"D�s�wN�\4_��
|$�]��V���`�KCvz�MەD+X�%�&�>�9%2�T|�ͷ٬N�U ���nf�r��u�����0!��(��Z�.M�hP���Ѕ��Zi��8	C[o��WC�h���j�t;��5��.�@�s�z߮|Vގ56t���+�>*��Yp���L+0G��%���� G��9�|f{W�a���Te�S��K�?N�`���>]���$�s���ZPۆ1 ���:Ж54�$�Bm�zS��(:<Y�}�wed����ȡ����E�AI�}��,sE��R4���y}���zcar�\`4H	d���ؑ���DC��HN����D�R�W?	e=t�̹�8���'��w,(|��G�s��y��w��ЌN|m�3HL8r�>�ylG�������H�o���d��GL��nAcD�(������J.#���=�(���� �	�R��y�-3Uh�V�۩�k�t�A��2���jc'z<h�w�s������{pM������POs����MT��u?d�%A#.����T���o8��|�<4Vʇ86���mֳ��F����R���1Z	P�!=��(}�V�,�Q#�)��|5tս�SHP]���3��/6���ՂO��)�*P�QN�r�O1�n���Cbh/�p�(y�c��$��G�r�%�ͬ�R/�qA�G�e�tˏ��8�\�E�]?��靜��_o�hFkB���3�׆�D�6��ĺJ�QjQJb8y%;nsv� ��L	m4\�^�Јؒd��r�>�PbEgvO3߳M���~�ܸ� R>�t����@\������P���K�/��z���AKl"�`-���j;64fi$�"wA�s9������+�1y���W9�V�S6��I��J���O����a��x�Q��U��F��Q���'��oȰ�9��^�y��cp�*��7?_�?Uܩ����Ǟ1�؞��hw��t��`.���ͧ�&f�}y_wjsg ӓغU��� ���m ��L&���p�X��Q����R2����|��d�K�QVԻ}��rLj�F fߐ��ZѩN/��4���D8ȩ�M�K�d�?�cm`A��GO/�����,��uN��r�]r
(t�|5���K��z1�������X�jg��:y��yr�
o,م���w_5����mҊ꣊������ħY�D��N�{��śym��װ{�O)�(�T��~���^�x�t������c��Ab�X��H{+�Ɗ���
�-� �L�h��e野�I3����(,�mC����:��B� �[X�i���H��� ��5Za[?^1��a�U�&��e��/NLY9`�X{�+D�<!�:����E�1!�/���",��n�T;��J��*F��և�h�c���Ѩ�)b45��?��BƆqJ@�Y����Q��� �����f������F#	���Ǻm>�w(�% �_�."��]�
�U�Ϲ}ҧDW�Gf-BU�Y0�yT/1�V�ާ^n��$!.O��vF�ma����w��Y����l]$k��L�
M����45�\���3y@W]�'ܚ�
;�N��C)�Z�i��6�ay�lz��Y-x똎�2[̪��G�[A��T��>�4������g�~��s�uYy�N8����'�W*䪧�Xt��w%�\�g�H��`+@{S��g5� �������V�mٙPџD��ׁ'GopL��d�9L�	�F�	���a*���5�J������Ҧ6��Șt�)�3�T�r���-d�4���v#�(к��>�ر���#�L��v'�t�Ǆ�VC;왒�WB�Ͷ�DѽTz܇ݴ�D�C4a&��%����LV[e2a��R
J,��ו���Kr��0�7�߻���⚊>�~�\5�-���f(��oG�&�ڏv�W]��S�?
/ו��!���=�ǥ�:~L�7��W��U�/���He���(�!�E��h_��GA�u�ˀд����1F= ��a�>�U�L��y��8v��ՑGZ|�"��h�vh�WW$�2�K ?�)�R
��J�k*������: �	o���WVa�����x:��!��Z)ϔ��D�x��}y�������6^�`�+c썍)���3_SϬ;��eh�3���
��]G�Ȅ�֞�,��h¹���*$�ɹ\f�c���W���<�S�@7���o�H��Msu!�c�JZ��b�AV���73�xN��pe��;����	!�G�3ٷ0I�at=M��0y@���m?�Bl��%�bk���']u�mV췍��n�BX��l����6�3��%!0A-D�B��*���s9��@�l�=7	45��_��0r�T��?1��f-�
|�sj�؍`�el�Y�f���Y��%A�i��%<�C���6M��)�9I�t����Z6(+�Y��A��>�۽lm�	�F�-���lr�d*GXD�����HW)�C*	�YðC\�j���3�)"������X��},)Kp�yl��Gx�T�R��t�_�)<��fI�G�Ur��߰��ۊt"��f�%���Jc�����I �i��X��śY�!�2���]h?�Q��/������GR%�q���s[Ix�|����UkS���1���!�Y_�g"��jWQ��L����Ɂ��o]qaW���vo�߁i*��<�o�	V���Eꌠ�����������;�Ɍ�v�4�i4.l~O�ߍ��H��t3'�>RsH� �b�0�i��/���A�-�Ո��T�>��]ſ�Y�O�00�
S�i��1��r1�m?U};q���@�}}~���p�$0��G7��r�\�����h
 W��W`P��ݞ��%�)���}o����k�?���J4<�y^��@���Hq*���zs�p~��'��_a98�����G��t� =Śrwȥ-@U�To_\��oL��8��w��Ttr���#�6B��YCK��)	�3���0��T��X�H��z���w��h�:կUؤ&�⌊�.zoY!Ꟑxe��
,�L5^_���6t<5D����r����@�]���Z��U�h  �W*��f)���������c�.<�dL'ç��0	aXP�|}v�����S�q����@�/
�1���Իe��/
}�Qb�h!��o&��!JM�GimS�{����M��}�8�t�TnG���`*�����d�s�*�32�R�ƹ-gҪh՟qJ��>�z2�"�q;�4{ ��EƳ��"d^�i�xƔ�T�X��l�;,n=ߊp��Z�u�
��|�F/��⏚0�����'��@Q�|k�eU�CR� 	ʱwY/�e��ſ
8W�����[C�Y��M��p
0�Ղ�B��ӥ4�
���I*g�KI@��Fːf�K��#냪I�j ƧҞږ<$��j�|��6Ͽ�<u���%|o|?;E�ByZ�֟X||e�G�AEK�6yX>V��8+0,M3��[�<
\ŗ��ᕆh(c�REǕ#�ܶ�TJ�T���ҤX��;�8p�2����Kc������ϴ��%r�h�(VЁL/f��/�
H�� �Jٜ]�V��R=q���<�l���a�v����r��[8��yd�z��8y5	�V�$0��`a��fC��`���w ];�hGy>�����4i�/f&q߃=`0�^!��P�L�H`q:���m����n�l��er��7��g��'M���^*�K��$�z/('f����?"�R���_���N�ڕ�[�1F���Q4�mݢ���V�i~�����1�����t6 ��䑄��Z����p�}g6^��L�{�(`"*_�p}ƺ���%֙���]�{O:��ªy2L:.�C�+�ܐ*:F���lRs^|�#�k�@1H�|{�2����]x&8��T(�Km��TP��!#K
3)[�sM���C��<�D�Xbe�C!����+�{c�"��:��8e���_nՂ��'[�.��j4�]�g��oR�KJ�n����تҁ�<e�J ��F��'&v���>�t+~6g؉>�1�w�y�FkeFrC���m��s�ۤ�=�3��;j���"n���i�q�9�[��[��B��S���m˷t�d*�f
YG�L�s����G��kacY>��f�J��V�ܛ�=�h^����3�S����D��=�.��a&���q���$o_@���T��scÁ�#o�"10rL���e?!_��������$�S�fǖFx�(����.аDk튊TA��R{� +������2����d�)���H�r�̽OK�1�T�J�0�%i�M4��T>Rhr���LEp��JY�Bh����r Y�ǬʻO�7����+ݫg��eM�Y!���ďaW�����AVV{�s?<K!R~�k��(���:޴�#)5����?A�����y{���P�/�����d�B�H񭈼��}��;�5��|����һ��%�"�$V~)�, ����A��3B���x�aސ�ڂ�ۦX$�$�3���i����d)�q�:Wit�
t,���u����`~�k��&N�>��'M[���NJ��h<s��Sf��o;����s*�mnD�<93��h�9�i��t�;�U�hE\�ͷK�&������2.�Y����2��#@�Mec�,[B�����kI�s���z���?r��� ����m�w�f�6�T��p�֓�H�qؿ�xt{��GVW��	wIE�)�S�Fm�ށ� YՎ-M,�C|F�������EKr;M��[M�y��Z��Q!���=J���A;������Q�iڌI�?�����"��D\[3��v	H	E^-����cq������ΑG��vkD�=��+|{�(~���yx{�N/�6a�/e�4�3FN0��tC��'#]^w�#��;��˲Z����b���������ïT��
{�b���4_�+\-q�	^��|M��`����ٺ�b���J�Dp��X�F�hq�'S�=Իw�,�iSW��]�D�[�?���E�D.όdC�b�Lα �$�JՒ0���'�n�i��D)���`�t9g�9�rh^���hD�G*�ޒ�)<?q9�)Y�8��@���}s3��LX@T�rQ�eC
y����	ꟲ4x��ɐ�({]��3�n�ڌ�v(�
H� ���o��pX�:��[5���h�����TO�po�tD ş
ҳ�����Y�hG/�k�R޳����o�	�R�UM_��%=b���Hs�"��Q��a�V����,�x�J/��	�NH��[��b=���\�a�s>#��,#�-�#*��̡"3�Q!kQ����<N���Q3P0]�oL~		���L�[��aa���@�R8��!���"�� I
��t$���ݠ������H���3�c��+r�ۼ���'��1x���F��]wz���n;(>���e����A�.kː�
**�U���2����sk�kj��>�⊦OY���v�T�d����e.Y�8Gh��D��7�Ö	���j;8�t�O��]^�%v�~xw�KO#�M),`>��	�_�R��X>�\`o9z��&N�k�9 =��z&:Ne��Ci��w"f\����#HR��\��&�e�U��{�6P�E�1b�É�`>��>@�N��Dx�%�񜋠V'F:�˜�v��M���ה�9'1x�X�{���{_�$=�rn@?ki]��*!�l��	V��'bԅ�fhH���$m��p�9�jf>e��	�HHU1!�N�}Va+��V��#�+sWjJK����Q!���D`\ �G�Q���;e�
��X�3b���W��b�����;(��RwY����{���۠4g���k*Ԇ�bXV��%{8�4�#��6d�Bϒ��$��	��֐� ����G���by�Hi�BX�,�p�h	���N���SwxA��u��Ss����p�q�U�ɦ�"/&׸99�u��8��d��$ox�q����8g� �a�2XqtMq�-��S4�i�Ɔ|��q����쥏���"H��b8��w����׵R6���3^�_fzEԆ�=r�y����s�x���rn�;�'���Y�#�6w0c�?TZ����)`�Lrv)���G�����)�L�j"�fh�?�mߤ��Ob"l+R��/�.R�'g�E�q-��i�g������_y"�	m����{��Q����iKԩ���F���Y�o��_	�Y���W�*R/W�i7�N} \9������y�͎ß}���t#J4e9$����F�&=���7����1�nі��Ł���uv��
��K�P�ы�Z\5�~uR#�kL)`�����/F���l�qn�� .�����`�zm�}�����t� ����A��P�n���K01��7�
?w�UbZ]�k�^�v]�ءH�+ �F����|��N�٧��[�-���Iq	��%�Ҏ*P0��~l@u����3d��G�@r�����B��� ި���)�Ko�mX&\
>�X�����۩�CU�����D�?>�yN�%�F���y�3G��^/���uV�VEG"�1ːjSʽGA�M�I�{�l�9��{���t�톁�t�Ο�a,. �L�0�vA�����`}B�K@�U�	�Rk� �((�dQv;�K�(A������,29�#��n�p��7�)�7a%�KnR+�D�.SFf�o�iH��F�b��>�p?��[�,��9��*���R����� -L����42H�������r���� ��a���@��X��YO����Mx�b���\���:Wb.�yR<�[x��;�W(���N�j>f�����D�'�B ��Q��߀0�G�WTμ��"ɣ2q�4�w3��D%�V�u�1l�����}Td��y�8i��7*-��E��V�ad����ǐ��C�9���1$k���kR�Q^f5Y����2 �c	�1ԑG?d#*d���v�b]W�|���zI��p��
�mX^ ���Z]4���-�s�|3a�ɍ���C�ݐ�����[^é�S�fQ/g.�����)Y�a�^���� �[�����T�ʋ�k�a�=�IY�(���u�^U��U�ϊ�Vۥ�����%�������0�9{5�)�;�v?`l�m��cUP+fP#*�a��Hnf�A4�G��k��40�|���R��y�Q�z�.wx	�)c�H
��w��!�=���A"b�r��#�=�
��=޷Q\U��R�k�[/ՍD�3*��4���'',�!%�s���Qb�F��3Wc�7�|7�gI̼�����~��-�����l�� �u<.e`���H��1?���ǲ�5�w���iw�>d�.�=o1s�{�c�]Ӕ����_��2K���xZ!��>������!��&�e��)��B���o&m{N�* mh��%9�òr�~��j(��s){[M��5���Q�P׺��WI���'�)�n{�#	O��y��ϣ�v!$�,��t����)S��[ѹ~��b~����Tx0ذ���^�C	A�ti+&�0މ��<��u2���Ĭ���Zx�`��Ʈ�ܹ���C�����Vi�i&��3~��|{]�w�u��,r���ǐg3��t�8�5Y���[�
II�x��v#��B�5`�ofU-o���Z�l�%��G��<�}R��vB��ɡ�X��^b�U� 0�0:5ݑ`�o&KG��d�詁�Cyܭ�L]<�8t��W� B�B�{[\�� ~d��]��x�T��n�䇡W�_	��+�����)G�H�|�4&���ϳ�%Ĉ.M�����U��=�ы7������1)�|�I�~�U �����K�Nv���6I��49@#� ����]jL ����-\)�WUs�Ggh-��RO^�+��f�8��]�>��kI�TB��w�{��(��/:��m��-��"u:�c�0횦Z��s-�<���
IR��{}#��{��i����Qsd�����bV�������|��q�1^��$�I���+���jm�o�Ȏ2�̏C�j��y�����N����_����.��,س�R�{&�)�(�����>�Q�U�D1{�)jǝaa���S�^L�͎\yYJ������<}k���sa`;ɸ
b�ɺ&6�l�*��z{�ķV^]��Wf����A@�C!�98I�`RN��>6L�����Ly�J=��;/�C�8X[8��kp
�G��%ܼ�Y[��m��p���,���7�7�y�3��ޭ���HQ�� ��O�S��E5M�����-w�\� jǊ�CQ�MD>��������FE��vE��u�0�"��a�K�5�6%��] ;[,�:�S�^-|���O�����d���|�
w��0 �D$�K|(߾@\���S���XN밻?�� �P���͢��ʤ
���� �>i�T��/7�,_������,��f�$k�EO�=���U�yV��3�<&���(i��Yw����B�����VUFИ!%8�B���go4��5�XJF��i6<E���F���
-�I��.Ƅ*#�Q��9�� 1�U �%�Z�-���-{L�C^���sW���_��m�<ė[�����rW�/��ˊ�c>�� ��,�6�A������t��Z2&�1n��Sη/e@��6�AVv���hS:��9Y�i��͌��s�?���v[=A��q�(�����LA��'�֥j���^��~`��.1w��;��B�vߗ�W����>��=f����/����,�_������H9����\���!$r,R�zG5�J������l"-Co���d���,% ;ꗅ���꾩��L@IW��YD8s{�Ji����ǇWaOIxR�,-�����:(p�s3u"�;�� I��tsJOL_����׺ķL4���ȑ3M�v	 ��������nZT�HqJ$l�7  �<�d�3�L��ЬH6�.��6A,.�~v�������O��od0T��\�%��/X�����m��J��p���.:�g��<8^aa��IԐC���;Hr��ZYS*+Z�~���^XW���"pW��ڛ���]g��ܤ��
:�Iw��Ӓr���c���g)�6w�gk+�s�C������y�Շ4�(�'EFQB]���`<�*��G2�a5�cD�o �wN&K!�O7�5��.�҆��/%2���=��ak�����x�t������|}��2�|�3u�O�)������s,�ۘ�~�X�۳19�#P?`�n��b���7���m*N���i��]@j��	5&f������:2<ȥs�Tr���pș�Wx�>�YC��:d���}>%{i�����.j���<�/��J�)������u�v�N�~�^�]>���Sv�LH�;��蝓]x���C���%V���ز�e�I+�&�$;'3�d�]z�;�5�3����,3�Ρ��7���L�J�����]�3�}CKǧ�������m3����7Q1��8�Lx�t,�x��zc��&
<��Hl�ۚN�dͰ���<5"��3f�;y�=2��ݩюs�v�Z�b;�aNU�xⅳ5��m��:��t��(���b���?\��� N%�fZA���<��<�d1�H�_8�&8���]�bFÛ_���W�0�ӹ�,��*�<���VL5��(�tq��}D+�9�����s�òb�Y��,���d[�o�'̼ء���vWb!�c˦�\Jl��mK4K�D�U'�y�~?�t�]���^G���r5�n�!R�A�U�VR@H9rg�CZ�[u�
7E�eȠ���cf�}!�Q�=�
�-����Oߓ����i�z��s�PR>��cV�"�x�
,�k��q�d���2�*�@b�ޗ���E�Y�/���8[��X�7������u���j�/��d��F���귕�+��8%�
e��k���2;"0bM�aG �TW�����}�����l��׎�{N?}j���M��;j^o�����{Qb.�)��*Z\��Ά_̽[\Q��a8�>΂���%<-B���~�k�%���H=m���L:�v�����\{�;���1�,t5��/c��G=�|ͤ�y�޶�f�x� S�ƺ\w��Q�K�,�`q3:�S�%N�J�Zd�÷�t79k׷=��|��'��S�Y��C.c5���}�&�������"����(�k���t'��ac+^Ά�C�{.;j~1�M��O��P�0٦mZ?�D��?�b�����}Q)PW#��s���H_�'�����K�?e2v#?k��-�������q�����2�?����:�D�B�9w��8�|-�ݞ �L,��Z��,s�x�Z��p�-(�_�c�
A�'ܢo��60&�m��Ǝ�b�b�*O�3��)��g[�5Ċ�bxƝӱX�y=��a���V]r�(��;T�0�������ٴ_x*~�!�n\o���	�!���o9��,A�b/S]���I �(�FRN�!FԶHئT_iW[�G�Lk��cc7��֏夅�}�Yc��*��|������5  !ޛŮF���4'�2略D\ހw@���Q���1ޝ�Q�DƄ�|����GxP��Z�#��$֬#
'w٩ 椗�?�Q�\���Fg�SȔ]\u�R^���)���khv�Qm��LY0G�,����6���b��p�q��2�SS��-]�+�p�F3��.;�yݛn_�&��쨍�����~�l�ʹ�n��!��*/�R_t�/�;����vA����t|b��Ih��՘��;����e{��0�n��|�_�~>4�J�; D�4�q��m��n��V�tY����d.Y��ȷL�T}��d%(�2��59^�K��x��&~H�b� ��6�h��'�?h�5�|r$�����m�T�]�fc@L
���e����A�^��Α��K��˯i���Xt�YMq2�>��q�L`Z�����b/� �JB�8>=
��d~�l`�װ4�ʣ-Y1<��
5��愕��7�K8������r�W�W.`��q��U�sG��l�2�9f}�y�"( t����#�
X��/<@����پ�$�w�q*چ����G��ϢD2���T=M"��[{`Mu�/=k�0��l�b�"`���/K|�qۺ�锅�]i{�qv:N{}��1pS�:�n?�����QjB_��7ØQ��ϕ(�R�e����������I\�+V�K����5���W��)UoO��(��L��Tt�R7���3� APZ���]ż�!G>���7�$����j@�.�v��Z��0/����Q�4�`�Y��Fk��ٗFU��*���vfIڟ(yLm���yû7R� uw<�����!d�Ny���|s�Wk��Gg�C��w��������H��E�n�V��E�@���!������蚙--}T�go�t��e��nb <����emu;O��/�����a���`zs5vJ�G��/��)l8�3)�A�{�����v�T���c��*O7�5�m��?/\�H�H27�s���j�19DQ���9�8鶏 �]��tP���1?�����]"r�M�q���ϟoA~�@�I�_�vx�t'�f���.Ji@i.�-��jºx�6IERd��ǉ����m����W��iǋ�A��?i n��-�D����M�!����"=� �y�����ƾ�0����
5���#-+���M���fx#Ur�ǝH��.������X��2�|��<S��l8`�T�gpI3��x��	��c�,��!_❝#��a��<HwBb�n�ɯ}M�+m��lW��4oߟ�;u)\4�U�ؙ�H&;�J~�䗆`�Tk��$Z!���	�2TΆs�ٙ�J�������0Ӹ�8�*|o�/�u�7È�����t"�H��SZf�X}�G��mѤ��r.#1��8U��{�v�<�u�U�䬧���)�
��a�z�5�xt�5k|�X�#/��S�CC@3{�s8c���,@���ǁ��
�Y@E&���MK�& 4f��n̤�A��Z����#���m?9�ɂ"���)��t��[�6[�W��K�M�qg�����	O���J\��<ܫH�eK�QS<-7y�1c�~{�d������sl���d�{aC�Ѯ"uJ�i5x"�����;�� �HO�
ksZ�G����k��"����_^{���
M>��B�֕��T����D^c R�$��Y���Ԇ8HȶW�$jn(�����hnjy��\�^�yc����/�y�~n��N���"�kw�H]��G�q�� Ĩ�)l�W{-l�|�?7�����]|tG���&�%&���@	1�pMlu�-�~Nr��G�獐���ͅ��á�Nj#Xt{˻��KCW���B�w�#��Ax�(��[�2���g���-J�.�JF9J{��l������
�I�+�����o�p�I˻�pg`烩	v����M��&��Z[��e!�����V���`L�v�VW�6ө�e�.��N_����N�b�٭�0��Qw�}���`��/�`?ޯ\�q�C�ZT#Vk&;����g�aR��<��`��p�<�wN���@D$���)|vż�}��
���7C+s���a���5��wk�ȅ)��V����<a)�O����f�H�Һ���R��z��+��9M�j�C�<�VlT��_(<�	��-Es8������.�*@�6����_�����0hU;�;uT>��V�y->���ƀ�^(���:3>ۛ�C�A�L���.��NL.U	�\�u V�;c]�R\u��l�F"�	��
��1Ko�U�Fd��}eZp�l���m�Qv���|k�ָ�0��Y��-?�"�a�M����'����*�Y�ԃ�R�n�o�8�2��P�T�'�H��;}��wvqcG�F�_7_
�"�j�	.5X,3+�������a�Y�5�z�]Wm+�H�H��D|�詨ϐ���ү@��#,�3Ły���M8����RHS4-���Ch΀���7�Mg��~g���eL�iS�1 �q�b���5�d/�hX~!dZ��Y܄�K�n�w�����\`v\����Т)���=C��g_q�]��[MI��mPFc��yv7�-�D�U�g�n"H�������!b�b��9(�Z�k�jg��t|�f����R�ޞ1f&��/ ��q.�$sB�L��"���	�j��_����(}�j3V:�2ָ�i�Nl��Z���U�o�ȩ����꙳|/mw�SJ����3�H곱���|�܏JN~5,�o2�w0/��*���^:��`i��A���_��9��W�J���kXtRQ��(���^����)��^��%�'��R@s}N9Ҧ�*�7%Q����J��h��-�c����^�C�bS�� �Q�f��ϩͣ��3W;��6Wڡ��+g�y��$t��(�z53���6�;����z%����[M�u�X+��U�!ᾝ��X���� �ɢ�D�����њ�֍{.����K"�Gg^���ܲ9��Ay�������R��a���� ��sH�wU?����^��0�W�`-�Zx!K?��
ڞ&�(q��H"EM/��))Tk�:�!����N��:%M�7q�x�[l��@�5�-�������Ii`���z���O��D�X�,��K5�,\��Q`{5�W�$�`�5>�����<j�����E�9��T�&ߗ�?��me��h���n�zΒU7�ڶ2�֨N�K�:�@�ć���x8��{J�g�WK�&����E�/D�����PQ���FE�x��["�ҋ�hߎs��w 7���CG�*Bm͝��Wh���왪�)���x`~�i�e�����|qې͘�W�h�`�α'� �p��0�^L���2�	���h����k8Nu���뇏�[8?b(;���p@��$2�5t؈�yat���םR�v�^쑊��JIg����X���%���6/ͅ�s�H�?��R߽x�'l��G��o�=;���N��c��_yl�{����Y@�1�~`^:�)�q�A����?=�#���f{r�	w�4�	�S��I�ŸO�O&�&0�J?��Pw�l��*4�Āɯ��syT�~;��w���6��Y4ʢ-��Pu/^Xp��E8�4w[�^
�YK�̣��8ط[,A%��h�z�}��!7���^��,<�y�9�<��N��FB���^��ލpF�a5��}_��ӣ���3ʡ�߀@B��8�'G��|���;`�{��;�X>��ݕC�h����$�j/�u���m~7�]uMe+y���O�	�r֞W>��)5_�x�%#/��[�R����3`���d�^`��)w�:��;�6	/-h}X�J���[�2���wy�ð@�],N}#4 �y8��)����luݯ���Y�.���,��[$	�8h�ebV������t� ��)<�Rp���9Vʘ�c�G��K1�:���Y��ݢ'���y_l\5{b��z�>h4

yz�Myx���lle�홲W��`�S7=�wl�Q4���$-�;
�7�f��T��&qJ7�ҙ�������\ٗ�/��s�7���" �f�6E���d�N�+�������aF8i�IN��aaP����n&-]��ԅ�^�
,������+���\d�:S\�T �����`Iq��;P����l��rIk�˅�儭��ǗE��;�U,��BT��x����������G�|�I�-�y$�C^2�c<����*�Ŧ��yW����4B���j�bX����%9�PF��{�9����3Y���s͘w�4!�z�������&�xʎ� �ۓ��>��F����n��Y��i� ��n���	7����8��e���v�$M�"-GM]b��r%I���J['2;�v���!|�'w��}#�P�9.Y֡8�{��;�}�g�	�Q�p��v{Ր�� s�`����0]+���Ӥ�ޞ��9��oܝ�i%~h9N���2Ӳ)�Eu�:�Q�f���O����Y�=OT�B:����Q���X��WpŤy��W[��`�,���=�%��S�V�2��tf��I�7�+Wm\�l��ć��ê����_e�}�Q�Cb^X�1T>\ɚ>�u�ٸ�Q�K.��]������mA[��?�e��VmZ�zV��x]̛}����z`U>�S;�&�~9Ϗ˓����.����U��-� 2�W�hm<��qꂼ0G��-4d���9�����a*^���Ni���1���(�튼�ͱ	�mzl(�I@/}�[�3���o��CaH9�i�9HZ<�GPNE���iiߍ�Ϝ8��e|(˚e�X ��p��.�]@ib��q<*����H�T)�c�Ua�Um��5�8�":/D���cI3�1��SF-�����>wc���Q�l۹*���kD�*�<VҠ�J5c�i��l�B^�i&�-�n�[dY�Oͽ5�P&�bau���<f����n#��|.��N����������.3� y�כe"�X�U!�ț����_��R�i��6-�w����=f���X�,�)�,�� ��D�WԳ�F�Kq�K��"������3��9��82]Is:�:�.�I���
�B�N	���	�zT7���H�x���k]?��gT�CK�
���&�O�/�f\�V=�����1�D�+S�l������y(3��4fK`|NC\G�.�,r)]x��q,(��29��o��Nq�y8�� Zp<�r%'-�`��L����\{a�0��{�&�&���4L���W�${�@Hj�i�.zrR��-�k��汳�!^�ei�������h�'F�QR0��]@l#���uAGG'L_d��������,�"*��>/z^@>ٺ��7�������]s+�j�{;�Lf �b$��d���0
��.;� �<��;��~~G���u.���~���|���T9�L���կރ�����	��>-_+��j@�����=�OJ1_V/�.}e��y��,�F�b��7얆kB~�^�|}�4�֯�c	�>�n�����x��c��,��}$�d��sn	� ;L��*Y�H���V��d��MP�&�X��1�i�?^���˞�#s`�W�`k.#/��ϱ'�N��pE��`����z7$珄ɺ�8&���-"g��)���k9'ރ��J
�i�z��i�p�3b�`��n����&�QY�<�C�����^̮+&垉�8�/�"&,���#e�Z�/�e"��T�u�$�o)�6�Hr(�����p6�.F)"��!�>�5t��H7��\5��~���|9�$u�uIX����jY�t{�I�s����w�b���M����D��つ�
w�g��3����Qh���h=+��
�5O�"AI��y`r\j��#T���{o4A�?6Dy����&0g!n���fCSm�~
�p'�F����P������������/_��r(*���H&0�'�%��s�4Sb�ʆ�# EΆ�+�l�/X��O�}� �`RKf�����rb����-T�SG�v0�q�aIzJ'�=��̚h4p��)q}�����Y�Hh]�0<q������/<�.BA��X#�U�>+�� �y��f�}+�Jo��IX)�_���ωZ�\����ֳ�����<�&�/��|ݼbrϻA?J �L���6�u]4 ����Ozg�Q���w�#S�@�ө�Co#�*��l�,P�����Gz#$Q����DZ�� �E�Wns��0�]�}Լ���9hq�LD�h�4�,l	~>�� .�s�Bgڤ�I��NE`�S�$���=oM�OÃC��CKj��Sմ�.�x�{x#���[��
� (݅��:�̾F�#s�d|�\�h��V�{�5++�?�R<��o�{�c+U�b~әJ$Gc�s�`�qB�ك�u���o>=z�����O!T�v��T��O�_n�^9Ú;���W��B��n�������4�L�� [����z8�9�C��Y��C��2��iՖ�M�|��� C<����7���1�x���~��[a��w���If�Q�!��3v�[wNB�2R=�TU���"��ZY���V�!��-��5U��.k��L��G8o��Hȶ�N=�D.�]���Wp��Tp��q�IE����_�K�͓�Նq��o6�u��Z�)�o��,F�y%���8-S9b�&�wn�t!U^��H�!l��P�� 2�j���(����DJ�����u6�{s��)N�Ṅ�ゼ��\������;���X�il�A>��#��RBWf^d��l�%0��<��}2}���/��~�g��ɋ��j�_��h��Z~$���|��#}���_���t����e-f�pb��k ����s��j~�~? ��c�tX�#��K��@.Bz�|���\
��ó�4>����"�Q��]���}A�q���@q����#���{�+�QN6�M&�HNS��|��I�{b��fIs��R��W*�չ�͖߰�ڽ#��x\./	'�C����?�m*)Gg��D���Ήln&��- 7\�����A
<=:ψ%gA�SBI�m=:�fxZu�����f	4v��G��Rk�[F��N�&��_����u� q����5zMN����\W9��ܕ` I3�����_܀M\�m��?��3u�|�L��U*\�zQ�e92`��	ݎ;�����-y�qd<�|QN���9�7UF��2����Xl�`ؗ4ǀ�%�O���O�6�n���� � B>��ϑ����p3��?�XL$�L�N�67T��fc������Ĕ�Xq4�S-�{-�Al�qP(�yL�fd��,��V�w�ZS8{Y�������n�Y�Y��0��A��K�)�K�z(A���ŉ�����g�!�X�s*6��2�J2���/�}�*8�S�o
�_��a��C�"ߵu�x���s�df��/yZb9w�7,bA_n�KH�D�8ޘ����j0�/K�\�̃�ٔ%�o�@|+��x��p-�^�E�QX8���7�C��߂&<���&}�c��?U[�:Fw~�P�]��b��f�C����w&vH`�V��.�L���������oUI��J�>:鵀.����i͍�.���'��0��A�G�q@���y}�1�c⅓7G�����ļ����@��$`�`}/�7��l}���:�y����h��<$�<ړw������t)~��7����Z"v��0#j0Y�� Aʺ{6G�Br��{���O�$߶Q_"҃�9]L5�������)<zXM*���/.:l;�)�"(�\~��. AAZ�^�f�=��G�a��} �A�~��x�ƺ��|���Fc/~Q�&����|��}+}H�iF95�{0���T��S|%^Nbܟ6ದc��/�ß�B��/��)��k��Vt�l](%%���Ѻ��E�b̵(���
n�s���M&���=��8ꤞґ�Xskj�R4.��F_��������L��(�����f`��I��hA�E����?��Ҕr~�ꂕ_��Zc�͎�7^7��� B��v/��I˹:@��N��m��]���I�<����V�X�Z�BBO��xّ�Hz������7���	G���j�p�s����(S�++m�Fb�F���)^���qj!�v/�`rӌ��9���@���MƠ�&>4J&k�5����y^=U\���P�^�I�/���E`�̣6����&o�z88�	�w����*��f�6)z~�f��)�UK�2�C#Zݐ�](r�m#J���慔���Ġ;Ȏ1zU�1c� ��n�����@�4�ܒ���ߡ���"�e�FZ/�����p7^O�u���T{��zLDi���[��&L��x�$�'miqY��	%��1���q�a���,m�7��z��񒚒zk���~򢌅�F��#�_Q�f�^e���V���!Y�wG��jأk��p��.�W�js�$�����>�?�?l/3{���
����6G�[sU�ZWL �
�*\��B�nuQi�/	]�����4��.�|�8�J����2i�-�{+*����\� f�A�{�� �t]kr-&h�%�;csP��4���]#���7��K p�lMS���`��_n���{9ը�z�*�g�w�ؕJ2VO����l�Qy�@���	o0d�
y���單P��3K�Y�wZ��Z��8��;p�@ Z+O��9�R��T��ΆSז�OGc/uR)7��v.����Zj ˡ�MJF��`nAd3ŲE�ܔF<fa�*���Z��\n��'bm�Oq]�s�P�A�筢���`lI��Q(�A����2Ϫ��W��!k��Cܠ�/q�5qv���$[_�p]�v�j��ZHɧ�\aV�+§9��0�M��ic�$��8F*�1
���vh���M�4�p�D���d%eԩ���͘������O,��ʎ��]��LP5m�	 l���z��*���`]��qIȠ�v昜�u�l��t�".q�d����iyO�ȧ�����ޡ	����i�gƌ�39k�b.��촣��-�'��w������_F@3i_�9�K�╷gn4�D���m�6�S��������)�V�]�U�g곗�5v��3�C ʄ���2@�Q�n�Y�d�`��jna�,kC�8�/Rɮ��Reɨ�E��U�{�m��*t�����-p�O��b��<�~����
i�δ�xp���|MwS��x�h�(���Y畅�ʏ`�CZ5�x��2��0 g�hD�D`�_��������[���^�~�{�|תג���f�ݨ�(;�-st�`A��O���W����s��x��^��i+==��|?(�C��bM�T�C=E� v��_^e�]s����Ajk�VLT�%���8�w5MOl��C�Yn;/�����������E�N%=N� �1����i�rg*�2���sV�O�ٮ躻v���g��o	�AD�����*�yL���M+�z��r[�������r��Xz�҈2��	��s ��q�1�t�L�����~6]��MNz����օ!m�r^�'������˪9��L�\*�oh�*R�ANV��)���uGi%�c���K�Z�.�oT٨08�z�)W��-b]=�Ԭ�15�$'av�bvzi�lɎ�"ˑX������kǹ.�� [ݺA$v:̽eb�G��Y����.
b#X�eC�$:	���5fX���yf�����,�8��~� ��a}��2/ �5FIL�����`Ŭ@~v>��O/���W�F�f�M㚆61��c��Z���[`=RC�Y��`�Y�o-3f-�N:��d09�QWVd��o7`�rx�\v����:�MI�qi(z,�D����?Ś�;�@<� �F�Y�pP����҅�uh��n��0&���ߝ��8C܄��&.x�8~g�l9O�t,@��V��S��R�Y��_�7� �(��<.06�@��b`߰a��B/"�a�ut��깢ܯ���{��d��-���?K�<��7�~<:�O����8FQ������Ͼ;�-RH��w;��eA��.�h[{��.�)~�,([�Tx��<��L:���*&+V�Q�V��v*<+f���'�.�yE�����R����H�C�]���B�|oA�|�-+�Ip9���=��_eV��@��Sg�#��T���_�neQ�(�p_0K5��L������,�>��+�@T�IP�ڤ11�7��o@T4q	Ū<ܳ����Bg�;ly�o�����.콳�<6���T�nc:� hq��P����� dlC�/G�,y�B�k�*�Ĭ1ꇰ�L}�<�����[�\��i`�����E��[���+>������_h=rc��s���������t �!OO���Xi ѯ����"|Gx����M�a��m t�È�W$�x������__�V��_R+�HN�?�3Pj�Ӯ�m��E�Z|�U�T&����@�׷��SZ��Tv?���Z���h�C�r��jIE@�S�tuD���.�I!���[��񓵜�l0I\�>L'	D��g����wAis[�H��n�e4��8�������M�Ng���W�j\��vgt+ꪦض�%����r���7��6�^��Vi'�X���1~ȓ���^z�gZ�)��g�=R��RY�}:�܊p�qC:�d���%8�h�uJLlSd�F��/�B½$���u�alW��FJ��^$T�Lw?�y���ޱ/7E�����	zVS���Xw%�!kD�/h��/��f��۟���|]є�S�=�0��V�)F)>�'�~G��&�L��^zǀ����<��C���������>|W���T 7����q'�>w�ȹ�
��^�SI���8�+å�Y�!�zs2�:��B����nP�O�1�~����`����I��O�N��g_d��Z��T��ju�]yx��s��).��V6����o�cj)f%2�?�p"fG�Ѵ�̠�=L��!^Zd*ְ
��M<U��G�LR���Jw��J�/��&��w�(R~`�����pf`�Pj�#��H�����sc�����h �e�R����) D�w2��	r���ֱ����/ԝ޴���	�e��n�M�c)	��,���}ر�$+���S�L?C�<ЁԜ��.���=/�2I�:|��~�RW +�&.+Rl�Ҵ2o�ё_�yΩ�Y���A4>�%B���<�Q&��0�	��1i;����I�?&�x9��=� L Q�+������C�I5�C�v]r�F)�J����b��6�)��b���F��38��0�|�x�zt��Gp�z��Jds?X/U��F�&���#B_ŋ2��h{G��o$.K��Oo�V�Ss|��2W�vJ {��̖�%����o{M��z9���̑i��Y�LL�2�#Zi��ü�����j�2���j�ʾ��s=U
1��KJ�M��M-���?Ƞ3���d9�Y�ݟ����@�:�boC{�^��Qb������k�(���b�cN�S
q��3��7U+�2/3]7�b��&�m��H���u���U�7���r��J;��yE7Q�'��%���Z�` ���YV�䐥�ΆB����Y#���/O�iIJ��"���g)d�y��F��ɡJr�WFT&��^y�r���4�O��h5�bT�~~�KX݉��d:G�a*Þ!����U�[c���{j�bͯ�߃������E�D�Ϟ!/��=��dw�t���$��S[�nțIR�|�ʤϽ/2�M�{����]��Т��P�N��,M(�k�oz}�#�^ou��_�b|�L:N��.�޵>3�g�I�)��=���)k��������Y@z#zpO(����6����&�P�$�&|ƭ��伛�5�,�1�Yc�( �����C�Ѻ�E��O�<S�tI����9AS=8\����r.�au���(.����Ex:��,@��&��$��{�.
��Ff��P�Pe�[�E�<�i�#�;&nr��������;�6>�T_�fl���3�zW73�c�����<�D�;�KA���kF�'}��:m
o{#iKҤ����FT)��bD��gbh0(�Z>����#;u�x�N����
��� ߩ���y��驏r��C��c�)[�@ȼ�p�K���A맿�L@�ǜ��V6�'�hF�4�{RB��. �m:�8�����D���9��P��ݨ�5�ق� ��c�gIPi!���|[C߲�X��ዟ4*��YCЍF=� π�;��&s��Kd�]Ql���@�D;���mjX�= Z��&VP���J,�-5h!�A�x��&u�icS��u��2��3��
�#gW�����R�:�;�,���B�t�R7��{���~�l���0��
@,�;���qG�.���f��ǚ����t"&�XJ����I6�-e�qI��e�![�9߹C��q��cТvH�F%Ϸ�/�)CM
��e�9U�#��R}O��bTe�沮��׌u��]P��/J ν�\��E�cVε��V�.���m�~[��=��E����4O�^Ŋ 6���Q�C�AJ���#MC�����o%Y�kr����^:D:k������B#ۆ6˞���0�ŔE,�+�;���s��V:0K\-_XW�
�t��^`
j,Oc�����ߙmoq��dH�d<~
~��	���?�����^�6��/.	��q0�U���7'�1���y�c2��~d�he�w�94U$\� mU��R�ޓڒy� �QOܒg��[�,X.M�X%�-��yl��N��C��r�-n]{^�����r����j��d�:�!���Y��_�n8ꄑ�y/̑T~=��d����rb�v��f�IͶZ�|�7�c��*[��^��~�����o��(Bz(	�h?N%L����n
�c�mXձ�r���\��u�,qK� ڷ!=��nW���(X`s���_�[�ccO=��s#X��D&�yˆݙ���"[g�(K�<Y:ƚ}��UX9U�����RAv��}�\��	N����v�oo��˵� `Uu�i7тzof=.����q�:��X@�)~���1�L�)��`Ow���pr��N� ��3Q˒Қ�8�z��0C+)�&f�$3���95�������x�]6���ߣ]���ʍ��؅�cI�"��!e�# ʟ�G�d�,9��TJ�F�o�M̰�9{&��Aea�EOo�����n�����ϩBM�Rѩ۠�3oi�ã)����[��q����"�#H�/>E|d�[kN5�&�F�s"C����&���@� �	֧K��]�����c��1�:dt��=�&�V��=OX3ߴD�u"�j��>]E�\^�k�q��p ����AӔDaj�Ҟ�8u�#��۔x�]g���	�,�M�$\
�t���ړ����F��q]Z\3
�SzM��=F��	QW��-=*��s���#y����dv�(t��(���j��|�t!u��>����L@h��y�.C��s���o���8\(��N
z�79�a�"=�%�S�l��x/7QD]IG��[��?g3��DMhҘ[^ӛL/I�C�զSgq�j &(����Ț.�+n�@]��h�kIm4��Z&(��>��!��a�u&JF�����+��"�����V�����ԏV�6��#r�GE�R�Xx����J�[E�R���.�Nβ�:[X�g�0p�`�fo��{���䲜�ʷ��W���2eN��~�g5�/\'>���G�~�������r���y�f`f��n��T_����"�?�4\WMał��J�Χ��&�����;���zy�_��S{�>E��DYAGn���+��6ĲQ./�~=y��O5$�%�U��~W7���]F�(���|�U��NA ���tD4u�Ի<��uԯﲁ�^.��1o��
?���{M�h��^j�[�\�A#�z>�K<r����q9P��=������t��N0*>l"��.���kUM��f����Ϲ��$���N���]���/h!p3�Reo�1��@��ccwd2�/]��F��I���<K��t��x/����u`Y��H3��k��n�0���i�����;�pu��q��_fj������>��%Hy�5߸���&���������?0��Vr*tS��_�U���K�yt�Fh<�780�T�d��GzGP&�o��K��w����F#dh��g3x�6���D�]B��(�Q��K#U������|�A�F��*e&=n�R���.	�$w:��2bshK@���߲�S����B`���P���q��S�XynPJ)��e�;*(���U�o*�������{���m`�{�L>E�:��PW(v�ސ�[�DY��N��_;�y�k�$ ��L�/�<XC�̓¡%����Q�$[P4#u��S3��4�9�#rR���*��Ҡ3�wS�hK�o��]������E���L�ݏ 6�g_���ØҌ�,FM��
� �z����>g���Z���Q���L��:4�$��v��Yi����Zz� з����-�՜*@W���|D�Ə����0nn�1��ߌ���kԴ�t9���i:Ƚ�"}o:�Eٶk+|���N|A�L�K�r/.n^�Y7�)�V����Vyc=C����[I64|��k�u,:^LH�`h��2�q���������w�ӹ��$�u�`~���|�Tdd�.�o��D1
����Y�kh.��oMk��3����rtE������R��-ů,���0i��+z�@@8��mic�x��v����&��$E�瑩���y�f��|{�����o��ZO-r�I�����	�Ƣ_>N3��J�ޕ������![�A�D)�dy��.5.�,�7��ޣ?���c���2�9^-<ո���j��EZڽ�w�������w�ԟ`1�4��T�/��6�J��?����b5s�{�lh%ֹ���͇|\�)��I�+8~���>�^;��,����@��^��a���LC��?/A���,��@Bj���_�Ը�;2a���ǜs�OG48޵� w���ķ,>s[x�5+�)^��W�a��>��(�x@����]�P��iAw�K�2�������^�oi R_Hs�Bk�$�9]T��X,&N�@=%RL��(����>r_C�$�0�̖�*�>'{��K	��b	�J�#���bC�V")�!���\i��)��S �_�З(o�0�]�Y�5h���l��b���:��{�z�)R����-�F֐���BR��Q��j��%��Y�:y��$��ꄙ=��b�(>f�W�ɼ�y��ay�u>��N�@L ?��.3��a�o�A�k�x��=:�-U����r# �B��)�?�ǩ�����K�~��X+4p��A��I�gh�-���*s	������|��(��%�<F�'���N���k�u)��C� ,]��XU�j��6�]��&Q��9H�w�vA8�w���WӯG~ǐ.���	 ס�>����p��uI�?��mQ 82:I.t;λo��wy��\7��e������uDnĲ���=���֦������/tp�@վQ��e��o̦�,*b�ˇeI�!��8�NJv���9'٣�E�+@O�������|6XF�_f���]MK3Ԏ퍟+�����"�����P�=��R���
/�q UN�u&ê?�6i�5�{�T��I���O���	��St�%�ݹ��n~0���1�]��츹M�|��������Ag�6,�*!?,D�g��>7��-�ذ��Y�و��2ol�d�'OY������O;��AVy�Do���[/�4�]�ݶ���R�n�-���GR>�M�؆S9��a�N��ajZ�h�+/]o.��^T��WLSDf�^���|C�e� 1F:��=����߄��xe��[���� `�ÓZ�r���r| �u���a��+�?���n����w��-�)����c��䬸D�,|�(78ُ�s?DDE7x/B+8�N[��q���Њx��~�_wj�X�g(M`�r�&*��/��WU	Q�=Q�7�a^�c��F�kIP�ۇm�3��{� �{�3��$>���0�����I���tA\|L�9,%��췬0J!'I��7���*��$.��z�O6�������. �� Q�l���?\�BW(�&�~tk�G_���d|�t�Tx�_�	�܌?=�@�G�W���"���1���Rc
���C�1�Գ{���.��g�O������Tq�R���>��i��f�W1.nv�`͏�}��x�u���O䎐k�c�0M�X�0Zh�M��1��k�}Ey��@����Э�2	߫2��u�98,�,��%�; ��tW	xooJ�S�=:��B�)�+68C+�Lj��|����Cbt;��a�f�g�^��W�y7M���~V���^'�cLM XbF��>ұ;�ֳ�-�Ob��I+��H��E�W��<��@���Q"���(��5��� ��xd��|t/c��jpf]�Nq�:$�团S!��� �������i� �,t}ݐ�|�''�S@���ҭ���~��-L?d��^�OE՘&��b��o/�~��l2���c���gyuggI��ib]� �(��Om��w�u��a٘�u�X=�eZ9#g���?n|����t��,y�hm�N�h�Œ+�� v.�%�6d1h�j %�����aA�̋B���WĴ��/�s}��R�r��i/���M#]޵���̳��W5��M٢Cw�/����F)�[5�uk����M&;\��mD!�|�)~�Z�i�8t8�~���^(��x��I�m6=&z~8MG*Ҽ y얘�]쫱pZf(R�S'�9��1�µ6��`l��5�&��I��]#�ݺIj�H��J�O:3u���b��.�Y��G�;�S���wm�vw�ѕb�h$�@�놼I�ַ�����@K��{:~>�����/�N�g��Z{62�н*�D,��U!T��ɯ�g�t���&��!�����;��q�C��L����d���ޔ;�)��T�A���v�3Z�dؿ1��Î�4�Qƫ=��Eq����H�
8���(��z�)";|��wh-:."l�u#��jV�,�,Ha��̬���3�C���u���V�u���f�.� "LWo��8�$���-8���C3Gz"#�K��2c���iy�=�	i��p��#�*5V*��$�B8��Dt�Z3��%w��O���S���og,f�?))�����@g|��bk���G�T�Hm������$��c�:y;=	St7���(zT����/�1q�%��#��P�L;��Ր�)8��d�_������R�.�į@�"��t���愋d�p�+���tg[���6f�x��1m��"22�d@?FwkLm�����i	D���+��tO�òåi������qxLS9���b���2�E�2i��0)�y����/��Rn��W�LKL�<�б�2s=>D��;���H��t��-@w;{��u�Zݬ��ƲȎ��h��l����q�^�;iX8�ڹW��&��6sl���P���K�|30ml:U�E���?i�K*����X`h7P�|�-@j�lxb:OF�!�5vC	g���`�]3xO����Qm�Q=v�/ t9�҇զ
t�qw������oF����.H�8���<�ҽ%[V����xu�����F�0���/��l-J�@�>Q.��_W�`�x�S;8���:$�����H)<W#� $�^�d���ɏ÷z׬ ��"�\=��:-����
kE�������sb�D��匞�p���V�-���x��!; ��~5�~@^+#�i�)\���4�M<I�I	��/�PRy��ۢY�pY��Ǉ�/�{���B�>�$�=� ��</�܄hI8y��i���e�)-�y��L�{4ubY���*�֊I-6�%�p�K!o�/��p!�~SLǛ{��ß�Q�m�e�dR-<��^�>P�k����"�<q9���z�S�2{��#�9��7���e�P%�3�A�V��hс]蕔�vo�r�>_�:pm%l�%Q�[n�1'�w}i��`��V�Ո(���V&�3��j�f�u�469o>�w�31cfK	F�\}�.ɡ�H+�ka��GվЉ����֧7���t5p���ɰ�&n�Y����%UX��P��қn����1�������(�j�0�@�=�a�Wө4$�B�!6��3en�o�B�r�Q ��p��C�q%�h�@���U.�N���V5�b�
څ�U7���ڎf��W���i������ �ZbBA����5DLn���������3���[� 5�t�Z,Ů]� vyͬ�<^�����T8�|��P|}j�I�[��Ӟ�8m��8���_	���*�q���4M�����bGDO��=%��o��3��:���6�1�u�E�^����8Y�۲�G�}����*r���IO]����kw�ے�P�������V;QW�M�,�8M�:^�4�L�2�	�ek:���]��2I�9�CpG�����!�/�Ԗ�w�t���։*�*��g�P���'���Eے�]�km)�6^P=N4�̶ҤT�g�P�s�j*�ӑ�YѶ`d�B�(�1�(��r�~a���ޮ�o���(�8����cKQ��C�34N{��2���f�@L_t&�*��a˹y%@�0<��&���Ō58C�ie@��	�G��H,�ZdX�%��t�h��x��	zô�j�GY~��;I[��#�t:�/�-��J"xag5�7�H̱.,|��E?�C��i�RO��F�%J�� ��52��B�v��zQ���\J���֠5nq ���|_܊(y�c
��M�������\��`���[��ɭ�ګ6�2\ 1X*�4��Wb���v�M�ӬboU~�_~<$	Qk�C}d��"p�5���R%J� �zj？wۚ�^���8�T������\��j���+�����%�~�3��=��K�J� �KN�-(k�x0�o���<?�k�y;�b�uD�@�%�r��5���Kʝ�]T1Nq�:��0��|����"8��������gs�l
���o�i��NLLJ򟄔
vwJ�jq�����S�X&.�g&v�ɠ}��W�s?�DN���}b�3��~���Ͽ-��Ƈ��~�iO"�K1�)��HQ}�we:�=/U�b�s=�_
-���(�S���S�ug�/$�
H��26j�Y"��A�h�#X`�J%Z�]�]�I�d<q�(��~�ֳ��(�㕴�Qa���C�7!�X�9c� C�VՖ���P=��-Bkz�"\��K����~����5v��6���@\�= Q��w/��H9K7��L,�-ifh���w(��Y��Y[��S����pp/6�U�Ι�H-�x��l
��3m��Д�MlŢu:�'��f}Mq�鰌*%���x� �M�++��r�W��/6���ǩ"�鿥�I����E��`����kx�_ď�\L�I�@G�3���e��`/i�</5$ҔFi��;��3��]��:ui7<������e�O�0�$���^����Fx��|�̰C��Ss��#��˼��\���K�#�IͿ���,c�m��<U��H����U�i?q����,d'_Շ�ɕ��;�,��Y��6��o"+N�$?�L�X�2�$$�ߡ<'���3���nb[�8��dӹX$�Z�C����smh���E�?1����a�4����7�2�o"�W���!�֗�S��s�7%%�3�N�Z5C��Q�M�ۻ���M!1~4X?����r"�ř��{�u�����	h���qjn�c.�6�Lf6��ij��`���2�@���d_�m�?���{�����1s����6t��a}~�:�^�I��s��S�9k��B�VA't�K�x�nј52�7�̡WzN&�	�$�9w�U�����ZI��fba ���E����zG��J�^�	pެH 7M����/tl�X+Z�0����x���K�K�{r����>O�1M,R��Ó(ۖ���]^X��p��ט���-l�;�F�,=�_7�5��'����6~e8�1��I���x?��%�W��[n��ϸ9���a�����->�E��΍Ĺ��/�����j��]Z��!�����BU��5��#`�;7�~��eХ��C��﯂i��=�0/��8�+hB�M���,\�^Zف���]`U?M�ծ�;"摱�;=�3�d��<�����G��>�>m���w����;���]�ӯ$�Н�;�2�[W�2��o�hڱ�ek6�h�3��yh+�p�&��G��KFP$��4duJP8��uVi�8�O����-Ǿ΂��0�H�U�yJ���)i�����16"`<�WU5�8N��IVp0���y~y4�2���� 	YN�����U�%��yg�^�w��.<��;��/v*,{ݹT�M������G�:�VZ��L�{����\d�0�g�Ow�r ��T�g[�����;���LQ�r��~Wj"�~�+>VΌ�/�(h+��q7�%�FR+��n�S[������4���?����}_�mfs��e�襻l2��2/4�6P��c��֨5ݪ���~��@A��T=��������U���i8�f�ǴQ/J�yΟ�$3ʖ#8x3X8�d���V{půV�rw�΀/F�W�[@��j���%�Y�Uѡ%��o�|�yL݀k�ԉ�ʚ<!�T�B)��+G��Ơ:��M�����r��q	"�y?�M�����a�s[�AZ�֒������ӗx	<��@$Q'�2�[)Ao�����tN�d��Q(&�<�;�;:�)*BYx��ڰ�r��՝�lv����������\v����S;�$ϒ�k���'�-�rPvr�"�~����3\_��{���YɷF���?k����T���[���0��`�?�`��r؟k��z���%���dmaY	_�WZ��ڼ�Q`����-\��ɮN�Xq�-�oc�Bk�x��D�@�r�:ôvoo*��fm�OB)X��_g��(_]W�����8����Q��-~�ɥ�������T<O�m�v�.��s	v�2Ts�nPU�Ѿ�dY<�+w|���Y����.h��O8��MI��q��/
 � d�f��>7�^*�j�ר�n ����Amr����"<P��ߞ�������ZW��^w(��[3z���;.��;*�܃T"�*f<�T�!�e��Cr�hJV&W��B��z�dZ��hG]����-|�۷d>c1}	~��X �'����V",�_8LB�5�m��U���Æ1��~�0���bc+�"�f������OɕW�.`}��f��Ugq��N�y�"�=�u��z�z�'��y����-�۹�&�è�׆l{�������9�b���Í���q�Z�vUxRNf��$�Ҫ[M��頌�`:��5n�-,�o)�.��1Z^�{�Ոj��qX{�.]kE�ay�=ߴ:���.wtoXH#e���Qʏ�V�E�B{��#��M?��ɚX����#j�D�E>�y �1�4ܙ��&VU�\��k3���\������pa�c!4c;Üf�߫s������s9RM=dP>�w�{(-~��К��l����g�,�(��\��m���@r%]�NAME;��G�4u\����V��9����:4A���B{���9I�jc^P3����&����=s���k�,�3�] �t�پY����G\��E~
Q���\���9�}�	��!UM�Ms)q_��S��A������@{z��_أi� JB��.*�k���?,�����(#-!oa1��'6��u5E�JoA�Y'Ӳ�+8@Ia���ϴ�7���3~!*��������ż�*�eX���eN���c�މX\�BU��\��ɸF�Q����ļkO�Z����A@��[�N�"$dZ�_����)d����X)���+ߵ~�����!��	ld�2�ۡ�25Mo��Y�L�煲���
��89Y�Q[��ʝY���$���]�I����8݃*�����L�c��Ȥ��l��ko}�[��~����!�^K8��ͺ7H�L�Nm)YR��U�+)+_U�=T�JSv,��|)�)$�i�pB��>�3�'7�9����Qdx�~�3C��v�r1n��l�I�����U���ΏX���JY-w�C�y�kku>\ʕ��y�e Z&�|���A�c��Y4B������Rf����-����Ʊ�}�t��&�8$k7*ak��>I)���e,h���.U��!9����6��_t�x,Vm_��0��9,ݬ$Tؓ����A~tL����+����\��3qL�d|D���ׯ�b�����ʇ�������H�4xK�ʵ�
ơ!m��}v�'9� x\۠ƠBfCF,<~˙2��v�����W�<96�}�:�L^p֧���v��9�m��ۜETq��U@�h諻��PE�ӣ�����c�Q�|�4���)�0G�{�jh�8K�q�m��2�Ս�[!�*��j/�u*B�ا�Z��Z~[���0���#�;M��ɆC�̼�S�lR�m��P����4�A!����'�t�A��e���q|hI�3>�L�5>�{@
���}�1ޥ�:|j.?p��p�D.Y[�ݳ�_[r~��y����Q��m�HQ]6�=�I��ʤ��y�G�x��lc��;>���%�����k��p���-��v:Y��(��>S�%�Q�YMM��W�"je+�+����fG���;����p��o�B�h�P%�k�j�h˭�Ծ�Y{w���!��>��J�[�l�E�?��CE��q��7: 2 -M��߰�P�&�1��RuK{j��I�M��B��Uc~�I]}���l���<��ώץH�d8��m����d|��H��3���1���0m�������U���8�ZY�xI�`���u������#��t:��]w���P�-B��G��4� lcVM�2So�ͼ*�����OS�^wG���V�>*k�e��13Qp�a��
�RR��a�,���a�W;���x6�K����2�՚���'�W�!�`>��;����ެ��-��0��{���Z����v6z��p;[�2�,>�㰗н���^�h� [ޫ?P�|(	���'+�GU ���� �QX�}����;�y�$*���HN��M;!w�;c�٧�C�+5-?4��7�r��REL�Ͻ�-�XU�O��
���[�kT;����v�08��Vׯ����c�Z����7eٓ����[�Q0|f9��%���7 _�s/0�o�|��b7�/oIGA3��o�!��yH��`��,���*�s �s�=��>(���v�$�DW����G�9�4��j2��V�(~U�F%Wq�S���OR�-�x�q7�5�Me�>��!�X�VǮ�ǐ/u~��v��>�*[�'Tv��U���B(�Ѭ�@���w�h`�gj�N��h�u��|�~��)`49�=G��>9G��<_u��do�������5D����\�$�p�����sV�a�ғ��!e���<n;�i:��I�z�p�!�v��iK+�u_�Uܿ��-¨d�V�>��>#�1's� ����Ẅ́&�f*�%vX.P\p'��u���0��?�L\Qڭ!դ��"b���X���8��8�'0�uJ[c�<U7���U],��d���oa��{U���N=X4�y���Y�@���5�E��y�ti��ꇘ��e%���6�r�3l#�=��<��,�8Y�X&�5�0���C�+)�|+�NP��9�%sO|q�k��R�2���˝�%#�m�A/�?7O��������r�{ʙ����Dp�M��i{�]Kc��M&�Ս��z��20�K<?�du�<��4����� �y�P�w, ��{=�)�}�����Hֆ�>�z�<�C�}���Yl"�����}����עF�og:��2?��L�T#�H:ܖȧS�$5P�\Ql�3|�x���	��V�#ݠ��V 	��8f=����
�-FȤ�O
�k��%��ID���ź��>Z���H��tOZ�̹(��<���oC�y[s�H b�����$�/�B�����X���K)�&+�H	_m=� _=bU���>�ʜ���>�c��T<���,���\��Y��y��,u���4��`��9�.]�N'���=�I\��mk u��06���a�����P<��HD+f��"�� m�D�]�.���᷍�����C�uҺ=Y1��kт5Qz
�=;z�C�#A}U9C�e��>�#��F�e����<ضlJN<Z����"���)!�iq�}��_��Wkʡ�t�Wo��L��m�Dʗ���H��?�&��n}�w�~?�&=lU���JH ��XO!K
Xs�1B��n֣��5�(�6�زM�rк�r�$+�ӆOB�O����R�d�2��2ZB�>�&7�&��-6$�U �g�8�p�����o2��J�x���`Wb�.f8&"֗cm����AE
���H��㥼uW̓�-^��G�6h�>��w��X+؏�t�m�~�i�h <���?�V@�D�ǀ֔��[��섲��R}M��:���$DVNㇹ؏զ�U�U�}O�p��I?O��!�`�+�:��������E��o��ȇ{;�ވ��0h�=��ɞW8�-=qI�<����4=B�'+6��+�YĶ=���Oͨ��J�-zР�!�|BY�!%#�4����{�Q�N^��ĕS)�x� 4�'��~��q�#�ӺlsYyd�����C:ve���{���/�F ����J\>�Ĵy�ķ���w��8��]C	���^�ޣ��aRG��B�>V4�b3Lj�T�,N�Rb�a%(@6��I��z�!�/��\��P�C
G��D��!�RP̛]d��u���Z^M��=���"41s���-L�������=��<��i�D�����"v����1�#k�-����5�P��s��ڊDs���ٗ�'cT�Fj�o��=�����1���
�a�Y6���WV��o�⣘�$��6��AV��?�$J�X3�$�l�%p��m`+>�3���� ���s.)mj]�f��n��
 ��� �*��2���7v��p��{!���09r�fv�]=��L�6g2`7^ӆ����4��䵪\�;�+�w{N6�a��ir��WN{�L�y�sH�e�ː��e߻���g=|I��J!x��F�,���@�!�B�_ǆ}�z%�n}����B ����u�I����Y�|x�{<�U�Zkl�&�D�&�/E��<%Y� �@�q_��,��ҺxI+��%�t���� ��V|�h�/CQМ�U6�u��V��L�$,� 6F9��1�>�@^���/�2���]���������F'���$�F}h���C_�P����|\_�i҉o��h\���s��zH����
c�0��}v�]��3�IԳ�g{ק��������ZF�p<ޡ����T��ǽ���nR&���
b�a����t���~K���mPo�ϳ�/{p�����&�ϐ�]gLf"�Bu�q;	�8�����1do!�=�X9^tB���nqoӀ����T��YG
������a%��W�uP$���	%���#�q9���Du]O`hbf/!��vU�{<,���J�L����s�f�뱗(�P4�"����2��u`��Xx���z�7��Eq ���ʡg�2�D3����$���;k���ɳ���F{KL|I�t�."�3DMᙃN)x �Y��x���U�S_�B]�)	���]JW6%J�'>H�rB`ۀ8/Q>�&�q
b:�K���T��WI�e���6��uS�Ȁ�NKqK(]�5o�-��鸃��4����I��i4�ԙĄ)�]61���b7��������Kqk���j��ʡ#�#�,���k�JГXW��'96� ������ѤxY��#0�a_X�vkD�PE�V`T��i�h�h}���L��aD�2�]t�M�9/tKjm��+�c8��S�x���1�F���SC
�9�z+ej�n�EQҝj�����
*��7������c@�~��T��W$lSX��	���=gotS���Wp4�x����.D��\48޴-�h�; ��L��*����xQqZq4*���Y��^ٿDB�8;t_��n�o;����m%���Mbnf����12�)����-g�Ui�n�g�_A�行��á�J��yd��	�Ĩ0S7,]����j�b��N2�xF1��ls�#�_��u��n�u�����x�5����^�����[��C�省��%��O>Y�ΥWd�g����s�[�Us4��)�<��u��c9Ox��.��v3�qs֚��UV� ���L��۩_%5��� �!�>]c֪T	�jQ�ϛ�3�A��x\Xi&��iSk���t�9��B��uv�G��"i�W�l��,xb����S���(��V�D?��O��l��"��үN	;��"������V~��mc�}�e~όb�\���l�N㰥2�Ur�G \0;]�F�f�!��Xy��H���+/{\������^�j���� !��[S�2��B�M�_�� ��)�7+W$iK�R�B��t����&��Ò��-���f��F: �z���0��/˕�,�3X�9�O*�pP1H���W�eX���1"���D�5χ�C�r�jd�V�+��m���x_W�RJ��L��} P���J����c�'Io	����sJॶ�	�?�&��K۪]��e7P!���Q���}q�f~T��ZX�C
"��e�4�V��$���v��!2̂�K�Լj�p<دj�qR~VJjl�>����&����������%78�4�Reo��Zbk�m�tS�y׏KSl�*U��M,�'�t�j�Vˀ'�����l#M��[x��� �_�Z\N��ȕ��wJ̧	h+d
;W;擝z�*�t+�χ<��&#�������JeW��V�eS⧸���$�b %I��]��`v�V�k��$�z`��<|�{�i𹞁�]����<6�A}:g��l�gw?�V�k�R�I.��n԰P��?�3;�}kq���v�]P�vD@5F��9��`��ҀJk��y�D�)���'� �	H���g֌��-L=7����A7IP�r]ڙ0��.w:��o��*�����H��y4��E\���l�,HX\o�[�� � ��9�P�/kG�H�nt�y�e������x}��WZq�!S�
Tn�ɓ�?_��;4�ob�]�2�'���g;<#��V
~�&�v[��t�3	Mw�:ӱ�9��-�
�L���a��-�m��[�^��a�A|�d�]�h�(�c�j�\��nch�to�h�>��9��Kmx�{I����A���=�vq<��r	��pjP@�ֻ�䀒I�������ޮ���t6�V�޹qF�2ܷ�)��C��k��+A֜�I�M
�y۰u^�bX*�yFB��-[�W�*�T]�2ʆqu3˞��D�;�t��o�Y�j������&N�0�>���e��RL�k8�pgdD3��Q�ÒXG.z�������.S$�}
� ��>���E��|ꪗ�\�d��R����ڽ�3 �ؗ#G��K�U)ُ�O�.xX�3X���2����z����#��/�V��-gyy�D�e�"V��+:Q��D�pȼNȄP�(n��EOk{8t�3&�K7e��7\�����i	����EEZM������<�3E،"Np�_;�t��)��QF�M�6\n�_*�yћk��99dFޓ9(<�Q�������Hّ�j败�1��BF��F��7�T��i��@;��[��)��
~m:�!�\�C`�\�Ö�G�!�$���(}����y�����[uN�$���XŞk��49)
A��ș�?ف�6|�E?xp��;��*|���}�;m&0�ق|<cW�^�	af�g.cfXٰ�B�D5?~@A����m�U}��ʪt��8-A�4�(Ȇ0�� ~u;*���!@��^����Q)��Q-@�"Q�r4��a�'3��_+������m���S�ji�W���%���h�ꌤ⾆�Rӏ��4�$nF�1��C�sL�"�����~�Cu�7��፩sh���oC����_�����/��F�Iǁ��_z��J���}h�  1�?��_Y�(�8����)[h�¦E*y�~6���]i[%m�P~:���t����d��1�Qr[�:-h���J�|n^�;�:���d����ar�����kTe���>_�@�-��y�<�V�D)u3Õ	f5����l��0�n5FH�=�����6>�99�K�s(�2�f���4�1�/�'�<HB�b�B�G�I��IB�cӿTk`��7N���������ө�9_�s��!m�{���H`��.r���T堻2�<��DҾ*�*�r�(�7�����f���
�(O�m��N�����?S���gmoA�����/�N���Fl�����5̓�>M`.qffsIm�+o�uMIU����vQ-!L�#D/klѾ~�3���Ѩ[m�MKY9u,�\>0�|��3��Zb��/=�r�T��-𝼵h�K`5BS��qe���U�ώI�f�PM�d���f_۹����a�X���m�70d�2�)	�:� M:~���`u�l��A]��DPD���m���K5�"n��Ŏ�!�U�*y���'}Z�(�NS��IQ�M��Υ�`o^��;���;V7^��u~~ `��"20������O�f��V�%(�x� ��� _$�Y�2~p>
Ͷ�tbՌ\�^�ы�-���`�<�����?|����ۓ�f��Z�;]�9[�+=E9�߰׫r�_<r�����{ <*�D�"pV��8�i���O�/��C���/H��[V��!��?���B]qv��o� .N�c���D�={AK]o3���M*u�'�+{Cb`���l�<��H-�U�p�F�����S���wG\�m�)����*~牗o�'��Uw=R��-Y͎�7�be��bt�:�e��$m�ԙ�����N���6q��C��4��S�6/#���;\�3��q%3x~�W�Sѱ ����g��G?W��=�y�}b�!�u�Af\b�M��E�!�bѰ�6q�F�iR��6���wd5
��?�M�	�Jq��Zr=jRٕ�V�s�ɉO\����. T-FA����.��ϩ�j��
(M'�~�)R��NG)�0s�pi&�Y�Q5 �E�[_f�!�w�N<����y�|n��Ǝϻ{>4���M�±�gG>�,5�9]��P�wϢ�X�);>���L^ݜU�r��A�����=n�s<�g���,�>!�Y�=z3�D���j��ee�I[�l�H(�����o��]�#�.����r{�����BS��pH>��[��>JY9���RS�HI�s�����}�����9a�x3��cƖX����/�s�i�l�Byψ��6�]��u��#qz�����M���-���<4t��l����Ȅ$�I�	�P�,��e'�H3�L���r�V��
Hm��O�Y+ߏ�`�a�Z���q MH� ��ꔚ�a�-?
��=>Ua��+T��o*��G{���ҡ�`��q8�5��g�����c @�Lʳ����ه�)��_My`�[:���ܴpB"	ĥ0�݃�'���︼�M�^�X�uĞ�����k���{N (Ӌ3?l\ѪXP���)�ry�~��^�SR�?̽�2ݢ��^?����*v9��n�Lg�\�R�5�Ж�@_u2��w����S�u�@�I�)ĥ�Y�~!����ß���S3E��b�j��Η����BB��e���8PT*0w�mqP0��3��#Z.��d>�R��#m�6<PC�x�Y�n3��?_*{����z�1A��W�i7)Vi�Y�ӟT�6�{<,{��V�JD\��(����,�u���c��7-]�q3���I�~[#�n�mq�S��}<2��!U��i��	->^�1"1�r�f+�Ep��lt�Qo���yi���=�M�{PS��Z&��{�{�o[���y�X��=95k֋�P��*YxH�Z[$�����VLA�"&#��%k�(\��V�c����E|:������*A���ѣ�ș������pƑZ����2���Ƴh�T\��Uy���5���g5�@)D��$]���_%�L�Gt	�ǁ@Z�����(a\_?pJx�6r�,���z�^��x�Y*lծi +T��Yd�ݛⰤ3�	�g��S�2C�RӰ*� �q�I{7�����X��_ �?����Z-��s��'nq���<���oD��½lL�2��϶r9d;)k0�Q#y��M��]���0,[�@���=�{��?Oj쥍���3t���5���Ve�2CT���8f��.撫:�fn*6���h���Cd��u�hgD��r�C�� ���,uJ�Y�6��- �%��{M��������=6m�
����?ğ@������2i��c�̞xU3*�cK9J��8��4t�B�>��#���vPRJ#.v���'D\��8Uj�V�� C��iW֜�j'����}f��O�&*Sr7�Ϧ��O�:�C�h�,a{�l@8a>|F��B���a}so�TG��6>�Us(j�C��U�M�zL|���ߑ݅��ɿDYv�]���ࣳ8~<�0""� c�4�h��8��9G]�4Ɛ|��vMY�A'��"\Opw��ڤV5,�l�|I���"Ƿ� �5_QD��6G�	�0+���]�]�����5f�=���:h�ݙEv�7I�	$-�l�)k9*��n5�ș�Noe�;-�R4Ϩ\���oU�6�o�h3���,|5����E��֮��90�7��2[o�x�K�ِ��໲2y��́���s���L�d����/)��wdSB��&�g`��y�L`cPb\*FCܲF�,r��sTH<#�L�<g��g��,Z�51�\J������,�w��|����+F��	dF�p?��"	G_�!�Y��N��wo���Y�v'j������3N��l@!Ge�z�5b�j�eP%��H��{o��ZT9WQ&N�����k��{,���g�˓V<+qH%k��rp]	����3�s��9��B��Z§'�	Yq1O�9��?�H�=.�ߚV�z�	퍀�;G���Ls�i���d��V�BܯЁ�!�H�R8Flkx�zp��5�fK�aQ�v_�]���C���LT�^�9:��y��9y�e,��ݎ��Un����4��7܈D'����db�������F"�wa�Eu`����4���hg.��1V=��[�"������0���<�����0`_�����y�/������ǝ���w\gD߫�c��x1CAӗE�=n�����&�9�b��`�x!�4N��G)*��><!I����]x(��c�����&۴+���q���T=���N�3�#��!a��@�hώ��!��[�4�<V�*6��m\E��@�i��Ԙ��S@ֺ�{�������. ��ˠ��^��
�Ƥ����7�@��HǤ�����hP�W�x�P�4f��P���(�0��B���a;`t�-3���UW�3��!ʅ<�5.�Mi����a�a�IJ�no�ޱâIk3���7��qABtac=ʴ��^}�t�{�^�FҜIR�-'>��#�k�q�Y_]`�ȉk��j�X�n8�l�f'�HG�� �`LĦ�Q�M+Mi�>�i���3<��F�E��x��I�UQ����R��wK���<������2V��q^��7�O�@=?5E:� o@,� �M
R�HI�ö��+?D׽7�}�%'�ޕr.�<)F�}:�s�Z�8�qS��P;[^d���^Z�m��	1mz|`�=�0ʎ1��2<s?*s�yk�^WN���bD߰�8�U���T�R�w��\?�^�N��s�����+t)Z���7�\*߆���y'k#���ҥ5���6z\�����`!����g�m�;���_o�yl:tH�{B0�s'�OLn`��o�w4[0��%�3�*$����>iAc��F����`�n�Bv{?Z�ȱ-�L�L�xp�Cӕ�*m��vaң��M n���$�%�D����\j"�qAu����%s����X(`�U6آ�>�&�<C>>��L<=��bAR*J6���,{|�B:��[��=���p�>\�Z��?�b�H�	������y����-Qv� P�X3q�0����OE'�`@�	=��T#4�JZ�"'p��V��"���H<��%BV�m�)�������D=ӏy�{��@Z/	�'��R�L����7k:=��7�y я�����g�Re���f������&I�x�f4�ض�ƒ��a/G1�=a�a��.����a����gӷ�������j�A��oa��k��]�&�H[�q�G��)]b��5R�|�4�ibf&T�l��|��{8賢���3���&���s>���{��5��Q癤D� Z҅��	���!��Č���� TP�ɃW�F^+E/_B+���U��"��WS,[���gWFį^�Jjs��`;)y��ʥ�Q�8	��Z��B}�)lR-�r᮸�/6r�<p�m�M�Ep$�a�jS�W�+�f�(��bYfA۬�~/{�;B��Zenn��E!��N�ܣHF��y�i�x�G�`���a(��N~M����_���c�-E����d��E��6����r5�[t)�&�S`�Ρ$����K���5��>pZ�h�jx
��Ga#�c��q�
(�s}�_n��_��L4������WK�� S&:��f6�D�������3����X�f�#?������F�������.�$ [	7G�"|��#^��T45`[#K�A��Þ��6����<�F�k9��D��e����j�k�&��*hv��CH�D#���2q����b\��9F	H7֔P�$��&��,ɤt�������R�yU�Mys���A/��V=�I����F�]4� z�_��/6�i�"+����P^�p�y ��F1�A�lZ\����[v���� E��uj�A	sLĳ��k㳳�Z�q�K���M��x!�v���q�I������qv VAT���]���D/�Zn���w�["ߺ�X�ؘ�<��k�+��=�������r#�?��>㐴mh�4�H3B�d�� C��5j�>�L �Gy�pq��7�AX�Y���M`)]u�l�aa��8t��j�°.����V��,)��m��;�?&��_�-GfR��Dm��Lؽ��g^
gD�Z��`�Z��/�i�9�t>D0��R��e1I��� t�$ǘV��;�h�mwe��hV\�z =�F�[#���E0i)��9��1{p�Az�5�fߝ2r�WUB�g�U)c���l�����
��S25�T_;;_�v����6��S#]������m$��iT|�>D�N�>,�V<[<΀.9�3��]�O�T3��9�4��zֵ�f�&�ݽ����<%�F��hLȐ��/�"u��ݴ�T�0����(K3V ��)�x�΁Y�7�l�+ �73��f��kC-��������w2��C�`�&:��/;۹~��������Tt{�7#�L3рF&�].qm�B!!�a��k��.����l���%�+�;��Q���7�1�^�L٫5J�+�
bG�J�5	����;a�I�+�c����E��Lʑ�JЭ	FXK��VMl��=��"9�{����'��o�<�����y�)�er�P���̻O$c/[�@{����?��ȶ@W�q�H�F6,�0(bIf�vd�CQ-�U�ŭd7I�M��������;YtG���|�Ru���^�.���۱~���#w�=�zG�W���"�-�d}�����3�D�,�r�y�&�"PŌ�f=������t5���.�T?f���ؒ��O��g*U�Ű��\;�Ŧ���qy��G�dR�I�P�����.�0�L�Zϓ�hO���N��T�Q���5w,N�1�����ؔ�Q���~ڃ��n�fK�c�g�6��k���i���������,�a�	9���G�-.KWRVaɅ��H6�Օv�@��&�M��q	��N���r�8��%D2��{"����������!@���R|��	�ND[Q;T㘱�Z����JD�;1Y�֐ 
���o�"�D�wV�b�kۧ��Q���b��ۅ�@�-�ܑe�X�%%w����������T%1�>�P_~&>j��@�M)��R��78��]���h.���3������K��2����p4��6�>��r�8��H KķhU݂A[�3�}���b���.���*����4��H�jQ���0U>O혪_BJ�17��V@�l�/1)�t_�*�c^j �Ba���,�
0���o�{����^��1TFy�,�R-~��o�lυ���o���}'�D�Ն���{aL}���+k>�ۘD�`��k��4���xeM�mH�����Dc�;-xm8�F�I�Bs��Sv}�_E�NX����
=JS-�8	�ˣ��Jy.[@�SV#�2��p�%��o��WC���u.����u�c�̄J�G�'�gu"��Yj���]RW��\�⹤.t6,���CTۄn�����X�UX+7����C��b��t�П��?��~+X��Ft�p�1C! DoY
ó�%ZM��W9۝����t����i6��2����b���B�2�i̛�jUK�=E�O�������	x�A��K��uT��N�H��f�t	�K9��t766� : �0�-�t^X�3�R]�N~ޗ�
/��OS�D[��v�H�ۂ��׽Qh�)��Ϻ�~��쑙:q�Vh�ݡ1���ev�	��5ޤ��Wg�M/���	�LnO�^
��ڊ��<Ұ�\������1�'�ϑ'd�`-�L��i͉PV��W5��KS�d^͡ԥ�X�^Z�X8��-�r-26�[3��Hw��s҃�����
K|��M����CKc�?�_�L�P������5���%����Y�T����߈�5���x�f��'<�����a�J�@���ݵ0tN�Lޣ�'�ķ��c{��0�d�C��,�3\g�6������\FTP�F\?un��&A}�`j�_�#N\����-������T�J��d{H'��)r��{������{_������ϾС���dL55�c
B�5wU�#����R�j���������u�G����*�{�������L�T$�5D����i���yAF���
����[�>�! ��/�=am��/�JmŢ6d�{��y�d��#�n��V��Ա2C-��������D(�b��~����g/�R��A��+�k{��٣�X=��5�������GܤB�w��;�	ٰ������N���5�R��wn����.x?A�̥(F'�����<��������G��tLò���C�}��Η*B�]���h#�c���i�=��e�����d��c��&!p�K6ߗ�F���%����s(�����_b7���fR����h��ķ�Ԫ�����>c�n���������"I+_�x�T`#ϣ���XDfHՖҴ|��Zmy�5+:Z҅��Vbk��v�ǉ<I����v�\�t鏚���M�b#=���b��7��U�jsT=��V5�TWt��j�s������ھ#�׺����J&K�yX%�*b�ݴ�k~��Z���C����
:KY���ǟ\Ƨa1���l�z8�j�
�h�c�^J��5��V��:c��>�m�IJ���ݏ����-j��TJF6t��*-Ƚ���\�e�(��$�$�F���"�'���-O�6�4�K�k��@����Y`/o'>��]���Xїf"e�_��`���xc|��A�q��8:����q5�:[�w|�lC�ǻ�@b�4�=�Yx�0�x�>t�Fw���޶"�����uCyL;���R:yc�u^{��?C���W7f� �sбa��������nSf��wҮ���I�)iߞ[��J�,�P���%�Qq��E<!����n���:��gr�b:�Ԯ�W���S�'HC<��;)k��.V��xQw��-c�~����V�;�"����)d�����o���W���K��\*��`��c�'�R[	[ZEsl��ny+kt�CN5��\���k\����6����~�짰}����a�-��$�,��Y oE*��91d}����m�\3�ڶTD1�((�d�
rg�ev���j
��W���'�/5ot�/;�CČ�Ӳ�F��T��������X�=7�/XH�ǁ�45r�v�m�\>JtR����t��b1e@��Yh�s(2tE��Z��L��[^:Ӕc��!���]`���#U�zë�?�M��B�4PQ(S�Ƥ/W� (q�� ��f\ަ���p���FKrd@-͍��/��wn�3F���z���6FG��e�}�--���+y9�����l�`�n^\����T��S�J"��A�6�2���|s-^z�0}/����
����[��(Y�-�@'Kj�'X�Q�qF*|[d�<�\��Y� ��d����!�Mi�g���ۣ�#D�m�5y�|�g�	�ά����c�L�f�GKi�U-�� ��NQ³M�d�b�U�- S�)/'���~��h�_������Y׫��I��I�0��@�x�k�X�����݌E�UW�7:y�����U���#L�{k+��=�_�t����w(�˩Bc�|�N�"ð��������ˀw��(jr�zHֆ��ڞ�CnjA�0��c�Fwkz#E�N��� �&L��JOz��G�H�ى�4��tWtYޮ���BJ�D�t5��~�k�%�?�W.�M�+cS߁�Ctڿ �2FVA����RY҂�\2^�NT��A͇}ZWq�X���Ih��?�����[0g�0rU+c �F��-0��"��G�����H��4N|H(�4�P��7��¾H�q�h�xjR��"�Q�6#�a�ja4�0�W��y���t��w�_��=Gm'蟧�]�a��2s�аEq��pѣ��Z� U`�T.�����C'��$���P?_M��#�U�P�n�D�P�,)�d�݌��z�ߚ0|:R1�`eO}�;��i���P(� 7O?A�bgw),�^������0��C�/6�-W���H���k�k5�YH��#%�����Gx�3V6�o���yg�/F�
�|��s���Km���U
c�\-��������p�ۛN�6z5�S3(�ͦ���;@R�ڴe���+xJnf�|k��TM#��~��Ii����s�
_N�4V8&�d��W�*�	����%�cc�w<���E%�jʿ���I�I!Y���su� �hi�5�c�"s"՝^)��˺.�ր�bFNi�d`a}�@��\��-�y���p	��z��3~['���ưq��}�꩷�G��f#c�W�Vp�3�r*����m�/-�7D����ܠn%� �c'�״�V
���@�Z�.Av�'k��A�d/p3C����q�����v��Le2��v]�N��F1"�X���w7�S��9��&���M�7�I[�����M��Ȍ��I��~
��ud� .B��||d!���A@ꮖ�车�V��׺�:�%Os�A�L����	� s��~1E��'-��R� i��Ze��XY�ܷƝ"�Żu	�ڜ����U=V�ݿ������K��Z����?�J݌%22/BJc�hA��Sѐ�w��QEr1�%�2��jn$�$䋦�x�z糗��<�7�9و��N�0d������i�H
Y/�`%e��o|��"q4��N��z�J�
E�>�C��iT��7�1�UN�[����C��ߒu���tj�%z�śU�3RmM�2&�дl��$悁jT�W��l��V�E�bJ��X�{Ci�ʺ�e�$a�šƢ�9)���J��턝��X��1@��g�!x�ֆ�H�h��Œ�ѡS/@���2ޭ<���@K����4��T��q�j~Ǔ�i�8�j��D���8:=�H�����s���l�w��b�Zz��'�;I����C��~�C�Sa����
�֣����h�@�h���" �%.Nd�9�S���v�V)�n��cq~��R�Qs���[f�D�<�_41���ר=2$+����'���W����_L�j/�%�BW˴��SV�R��Ђ�bOc�K�w+y�v�K�'4L����3����ѹ��$�lll��M�Эwܱ6��n[�����yXф�j�������p�n�ߢ�9ս:j�#Iᚮ���W��7:�A�Txijqh�ޮ��2�¡�ا��쑅�{1� "s�� ��;�Hķ�:����s�I�p/ldx5�� �Hp�8N}?yڟ�A�$(�?�E��H˦�Vջ��~~�A-��GAC���|̃	~���{��VA\Ul�|{� �ϲJN����a��T��2�w�՛�Zw��V�L�5�H>�y\7��s�˟�3b�8#�	$�زϳ��A���D2���6���k��0x�?A,�)SF!v�/���`�ؙ�	��w�Wb�pO1jE�!L�D��VY���/o5d�=N�n��W������Ka$�˭W�&H�b&�?�^�N"����=ea��g�И��%c��<ʋ��0��sNw���Z�tPO����Q11�E@��{�:~��:n��GI���T�Eǭ�C�U�J�ݹXaF�	��Bv�0���4�v>�-��V� ��4�r�������A� $��[�G��1uU� ��!�@(�0*%�q�ͦpA�ˉ,�[�~d�evA�x|M;Üк�j�(�3�T��2�]�!^�T�w`����D,g
"�'�Ŝy�a�͎K�S@O�9CNԠ=P%��ɳ��j$�9 c��Ic�^�[�4Kwr֯� �FѨg�����dK�8���وD��9��7������I�$+����	�9���A ��f_g��.�jӾ-n��h��^�p|�����~�e��%����[a(�+Jxx4(���u�عq������!i�-�9�3S��}4��X�8=P�����׊�#�z�d�R����)��p���ɪ��ܾo�c��+�o9a�U�[��R�M[�묞�:��r�Pp�5��D�����{�N~yA�z�6�Y��N�$S����d�����Z��L����u�d0��ʶ�:����Ge;��pԱ��$2Fe8p�v�_�*�T@!C�M�].Ӌ�g�l��\[�+h\�k^��*��X/EvNCP/1]�@?^�Mr�AH�]?X���@�G����.c�K���/)�S���g�������w��m1�����	�&�{ܦ:�� �n�ѩ��pX�8��v��2���x��pZ(��9�'ߕ�X�)����9�
�L*��m"W [;g��G���\�Xe�G?4R��8�0&�+I~©j��ֹ:��B&�m�;�����y�	�n�,�����+����f�G8�70s#$?������[�����>=����{��t&3���Mz8�*+��!@ZVz���Q����b&���\t���?�n+���ۢtkеL���<5���B|�Qڴ���{�:�٤H��Nq�J9�*w����_�Ah��妻�Q��x����q3�9i��e�Vڝ@q{[���Y�t�)��x��e���H���ہi�������P8�����ln��K�O$�T�s������ �6���n;��(�fR�"�I��[������3
]Ϗ~Jy�*��&e��q��}y#�����4�⿔�M�\��<ڍ��oZb�x^:��/�rO�IS�y��(���W���2;�䩩dL���_���0Fcݵ�c�s��34�)��H�~h+��^��@��ñ�*�e�M�Òj�����W��� 4�	l� ��� ���(�&J�ǧ��t�/�<����G
�
��3+����NI�kS-�Օ������3K]�a�U�k�g>G,˫W�fC1<�j�	��o��f�c?��!̷�vsE%3*S��CRv�����r�+꺸XM�<��Y��+n�j�����ٲZ��V���X�=<��4�Y� ��E6[|mH�S�㴕}�oZ����2�I̦�&e�D>?y����o�	��$5}�i��z�N#�>t�ev��g��v��~χ93�_�t!�4]�^�B��q��N���RA��O��|2�;(R9g厊K��N���M� ���E�.�qb�fU�P�>(��>�>?G捿�ic�N�ћ�v�c6ޯl\�/�h��/��]m)�S��iN�әsv}C?%��Sֈ����=�&�P9ʃ�L��wi�Jœ�	�U�<]�x���r뺸t~�w���4� E|�|������;�r������)zk0L�ӭS��U���00��śu�j-�h���m������<¨�!�s�C���Qj�'���y]���K��: +�AzSɢ�j���&UTFW�w�P�_1�zG!��>Dcp�ʛ�p��E���Q �H���8e�5e�XE�,#ix�ĥf�����M�՞d�~t����|��q�y�<3>hw��L'n��D9b!\�1�%�:�����7Ɍ��Ms#E�[a4gլ9�DC:A�3��m����u�K��t;s��&�����BM)L�J��z���l1u'ˢ�<�{�0w��m��_ Uiy����Ri������2��4����3f�C���_�+��	�8@D��F��T�Q,:�"�E��dt���?��S�y>�'�+!��6���L�&;� *��L|ҷ���;Pk�������H��gH���H;;�?���� ���#��/��������63�w�`��@�Hó.�� Y��Y�$�d+�ʉ��U��_C��}�X������:����-��l����j����,f��=��I|!�	+�+��ĭz�۶;C��~����`%`~�
�z�F�N{c���zU�Nn��!�M��7]�f����x����_�f�C�~��F�Լp�5I���~`*,ےB��ϻ�R���=vw��M��7w�F+uډ��������0\ᢩ�47�N(�'J�D˟:W-v�N�9�px�~���Y�CA�-����7�	~��&�I��k���q�+�m^��&��tX�7(�1"�����a�iz$
<��5J��1yK7�ytVz*��8l[+D:	L�˨�0>{�IZ_4�Q���9>@��G_�$�1�m�;ו��Vϖ�jԋ	4s`�i�~�hL� ��AꎕzѢC�6�|��.&L���g�} $��F�s�/S�\�;��t���y��]��\�rƙ�mSM8ƴ�[�/#�A,�`XVc�?=[k(�ބ��7ڠ��M)7OT�e{�,��i��=�
�}��#���l����H?z�h���+�cd�>���b�
���e'Z�ɔ�[��*L��s�Ze����MY�s�m<⮛w�`���m�������N�}?�O��֒��4�ҽ�3ŋ
-*���Ŋ�ؓ�¼�pU��R!�Y���葫g���e��la����o���#ġY�X��B]�3P,$k���r,	���B�3>V�?IN>��۱�>�a����v��m�9�l��,Vf�e�������+��}�ɷ���͔�=��{Y0'��:��i*$:v]����l�p�R�D�n`���H ����z���P����-��$� �E�?C��\�8�9���B���~��:�$�jp!��j��G�k$du�(� ���� ^�i�G���֏
��O�	J��Aju�<��|�����ܮs���(_<����LPm?�u��8�b�pu����ٿ�����u������[����{�Z 4D��]5��K��昻�$�������ቨ�/���u�G��,����:��~h*����nx��,�+��d��4#��:i��\mF{����]�3@ �-����ƽ�yT_�M��qކ8�])�6CV�x�0C(���"��
�VB��V��#�<a�E�5�����{%MQv���*��Aލ�E%�V{e.�Z�x��K��YIq�A�U�������*	��t�4k��B5 �=7b�3�JI�`��J��n���I&�Ќ� �e��2 ���Z�06�kq3�6^&Q�P��b[�L;b�uczw��0��̧�o�h�2P��)�P��
��F�NѾ���F�2�R�x)�	�bI��s�33�\�=�(�9��>f4?̺Ս�8����B�hKbW}_�����tXPp�1#�P����=^��q,FYBL���?�a(�����b_�my�n�G��������+�d�~%M[?�<\�����d��f��5�	+�N6B�[ �B#�̧���+��9�jC˰��6�P��9ægِ߿)�N����?,ͨ΋!_��"�᝜��8�ΰl�k]��,�h݁�s��\Pf����Y��Ma>nb���5��O�}0��\cZ���ٯ+r���P�����l'�%�}�}�"X̬�όÓ=ٔ�2��:�=8<��&�6���}�T�)���A�hd9f���,�[���� *ݾQ��Q.C_!OW�Z(K�B��ٽ��n�_���f#±���f�zjvö�J����4?'{��mH��Ȓc�B|wRJ��P$p<Jx}���&�#Ê�?��9��ozJ� f��/�i�%��a��09���k� ����PtoC�V���%(+���|@�)�kt�&�����c�b'4�^0W�ea���U!��3���9�v�%]S$N���6�Uu�ASe� x׬�F�8٪*;q<>T��3��1���U�CA#�ޖ�R%�O���t^�8An:�q�����������̐T7)���Jr9{�0!� ���杮|9���nB=��̧���-�y��y�ʬ|�����I$�a�@yt^��Y��;4Ĳ9���bf����e���Pp���.-��,� J�`}溋�8A�nTD�F*N'�^�cb�=�NI~i�I\2셃8��غ��6�]���`<7F\� jJ/ k0��ʀ���Zf�1Y�Q1F��`��7�s�����5�ǽ0���W�;41��9B�������k�[W��ڿA1�4M�VG,�۾��B~?2��S����㐣f�����3�W��@���B����x6�(��V���G��qH����*��:[���P���7�0@?��I7��}l��
���s�"M@�0��1fz��p<C�ȭ��L�.�ul(��	�]Ex6�|x[��\Fk�:\%H:�*���I�[)p �@ïS����G	?W��V܅.��J���Nj����Vo��}KDݧ,��O���ӕ��*�4�G)�)]���e�9�8�O���p��r���&�9��Z�<��B2�X�味�앲B��B��t+V
�ǂW�,������s=���7���dՄvyN��Ù�RT�0Ͷ�@-;�Ԑ�䮉"��<ݑ5ۇ\��y8�9��9�lGߜ��z���S���,�h��"���o=�l���^��~��ߔ�����'��-9!n��s�X[��LVv�����h��N%.�hw7�n�RG!�E���2�jܞ����,T�43Ar���&�C@Ѝ(�}�MϢY2���{�0��~P��7����~�����O�Z�w��{U�m�qzA�/�
�L:��D�@��љw���!����c�-�����j
�:ݱ���u�"��+��+��{
W��+x�מU4�6��w��/�k.JD.�xΠ� �E����*t�Nc-|����gc�1h�L���~��ݞ3R���$����_������`���Q�t'|Y6��R�˼�w!�����;|犿#�Xo����r��PZ�Xl��P���p���2@�2�:�	&�!@��NZ+�os��G�3�u�K�R�.	FM�5�UqgtE>FM�8����ҍڵH�(����u�y^9��^3��Xb�G��	�8[�k��8�I����N�劧���5�}-�N��8��pu��|�����JS,��T�%�g��t��j�	P��@����<�H���:�]�9Er�+��iRO����Tf��y_�|�%I\L_��4E��k�6�+s�+ִ�elN����2���>�w�KJ��X��r뚜�@G�]]�l����[�>NwۅeH71y*H�����EO2���w���A0���k��,ۣr�D�}�r#��¢�X]��%��زi�.ǐ*�u��eݕ�0pP�^����u�C�xv2�#ŐP�S�<�$����{�� W����ܚɊI^��%OD�:��iKlʞX/_���@Af /�	!�6t��s|l���QA�[;s�w�3����9��/�U+c�	�<��)�Q���e�&�#5|�na����5d���v� ��u8����Wj��T�3xa�G&ąm�s�t����՛wP��)H9���a�<������g+� ���CPլH���D�b��;���t'9�
[�>l��8N-�l��a������#����A%/��9�m��u�$��5{�����4�"���[>��$?�x�����iľ9�����@�O����H{# ����1�~�n _����T��⳱���������4�<؉2<��1���wS%5�i��N���V�ʛ�dr;�r�;�O����7�o���Ρú�㝊��.x[��r{g��zy�.����;r@ys�����b3Z���r�1����M!��m�Qc��dy6 ^�tFӅD	z�Ҕ��X��.�r|�54�%/�ͣ߱r����,��i�GW����l~@�BIt����D8I�� �������$�Q��� �♅�#ۛ�/Jn���6�o���c��=>�o��&tɸvV��)P�U�K*��������f~ �3�R����{�6 ��å��y�z���Ն'�������F�����|�Ǭ%��$$VH��|�|qRC�r���=��L4����r�#ڿRr��ϥ7A��xK����I�7]��#5��2΄�m�H��<rV+q�d�!~�t"�K?���?)�~����p?�f&�L>��A��2DYhr���{A��?h����@�k[�6�Jh&��PUr�=|�q�Pi+���ѭz!h����X�c�w0��_?��J]C�i�7YU;�>�Ę&�eY���T�b}T{�
\w8l��e���9�X3Q�TҀ=N�Ӝ=��h2#�y���/k�/�@����DՓ}*![�R�-3Ͳ0K%N�(�uoϏ�za`(�1���^�di��S;�'t��o��~V�?�w�VNtT��<��� ��F	vp��b��a��״Δ�;Gt{��SQ�d~ R�{ڍT[�=fv{M�
?O����q��T�i�Y6��$��ax��+��8�0�ULP@Hѯ�|�'7�V��P�^L������8�@�o Z��ݷ���)ew�f���_w��8R�X���n��qǔ���j�\��ǚ7��df���kK�C�.7�������I6u%~�0C���x/�?}b������dJ�������T����U��IT��'���W@ynd�,�"�7M�;M�Pϸ�3��u��T�ߞ�LX5 ~}6�����4C8���;���-��)*�����Cn"�Zhm�k���s[g��!�Fb�΀*����lP=R?Ў-�m����[%k���N�m-�+�ٓ�@{������YZL"�$nN��G`�w�v��8����gPy��bɥa'D�Q�cH������e+�yh^�W�����a޻�����s�ij�nVX��ѬZYp2���2�K�k"�w�|;�8�4k�/�a�m����H$��t�K���j �@ʏ��=`a��@Q���Exe���?�G:��#<��O�W�m`<�Gk2�z'�K��;L�kM��kN�k+�/sQ���)'���@W�����0
\
��$PGȏ�}H��uHO.�7g+`��Ȳ��2����?9����|{��6o"d팓��a�-5z���L��~'�\�����J�=��M�����Y�f�P��9�Yn��n*�$n����RB�Q�s�A:/yLVd�>	��wNP.�ʱ�ʟ
��x:fRT}Z�\QU*~��dM�n���5y<�8~^8�+���O�YY �d��E�:AbL�K�j�OvUd��Ut��n�0�iޥ��	U���:f�,UX��Ug@O7��q�C7R+}	K�`�f���{)\�?��N�_�C��5e��8���p�1�<O�,�e������Kw�a,���G�5�����Ҥ��*�M��l?mȴ�`�u�}�`�;��'���_�@�M͕ar��� �Y�P0�ug��![!�c��" �����ɵa�r�t����
�'߶�v�wǓ�[̓�Q�-bW����5BT'U��~Ҝ�<-Wca�����ʌ�O[@ZZ���u���ٸ=�4h�=��k��������;��� Ȅ��ބ�>�����k�2x?u���ǔV��S ;��-ʍ��>G%�̦8��vI<i{/.���
K����G�8`U&aE��_,�����]Q��O�x3f����0dF��5�g	P�H"~u|�k��^J�3��O.91�3�g����#U�
�e1<�U���)+���I9�R�z��}�AB��I�|(;E-�׋R���y���>�j��4��<�W 즻!�0� ����?x�]�>f!�Y ��ot^APW��
,���LĎ�K�s���������H�1��M8\[����660�(я�Lq���8���Hp0��Ղ�@!x=��X���p0�Yb-��Չ�a[���K���xn�\��"��Z��l,ύJ��O�
����CkYP?i�6�����r};�����̝������ Ȝ��V0T�h|C�F�"��GAinS��pzi�����^&�����+�dO��� �Ts�V��NQ���]���H8������me�О9��!���2��~?��0\���KB��(	�����5q�{W��\{�8�T�����ô#x����)��t
�J��h4ٗK�Y�;�*)�6�r��g��ɛ����9�M��� �!q%oJ~�B�E��Ժ|��oh<iʮ�#h䢤�/����޽&h!�����K�dy^W�/u�Rajj�#�O*��;�8}*�8�6Mv>�|^.�]�u���F�E-��9���Y�w �v)���Wwy�^
��d���	�آ�Y����Tz�����/\����-�o���W�[��s����3ѹ�ӊXe�������Q,�4���POw���+�E���ԿtJ���p�������~6.�<�Z<�� �.~�MuV�7e}�#�*���~EZ���}|s�_[��� o��!F�E�A|iop��A���#�֬b�iaVf���.�^��|�f��0/:�%� ��c�o���Q� ��zL��s`'��� �5���X(�,Okn�э\�S�&V`��|b ��4�i��	6��}xLAom�$������bJ�,̳O��%��֕D��ט����w�.��le���1�X���g�4- �ޚ�A�!�h� ޑ9��&�i0s�(�4���A��z��m���ڭ ���O<��F��e�^�����jP�9/�˃}�?[�����]ߒ�N����I!���%i�m���5��b�!����X�	Lfx�gE���ޜ��OVmw�m�_/1��c֝ek����X�]�>�]f�:����@�;눭���|�]�I2I�er1��;�F�\��[Fy���ǎ�� #�2�dC��khxÊ��L���*F���|�����&}��Dw��3βڕKx^���pCj��\e#�?��9F�t��	�y3X�<�G���y�^��m�q��A�.E�ڛ�90���SB��N�(�ԨL��2�Ay$iҷf9��|]SDs���^�ߢ�Gp�>��ߨ#�w�_�|9��ZeI�l@��uP���0���0A9<��q"���ތ[��S��#�!��!�N^2��qЃ=��_�3���h�7vk��7�P �����@����k��ɏ�3�ʧcI�u4�~H��J��f��:p��s;�C��y[�)���=>���1.	��(�
)4����y�������<4&����=���b�����"a@�����y�`X����O���q����N޷By�����h
�NL��"���z�����=�	��u!�K0X�W:/a��\оM��U�M�3ʭ�RUq~�7�v�\�}�W���%�[|a��%�
ƃ�ۊ-i �E��"��^��4�fEɶ�H0,���m�i@m�,����+:Ȓ�L�iScBg(>�f����3d�ճ�$�}��\��]�|�mJ�[,ǻ( �瞡�Cۗ/�A�	���~b��l�����d��;���ǌ�6S�jj��4yĶ�u�`}Y��/�~6��;���`BR��v����������EQC�W�0�&�J��hC!�ňMț3���y8wZ�y��zG!��)q?��G���%�e�Η3NӃ����C��<Q�[�V�)�li�@�k޸����M��4F`����v\����D�>A�(%Ê-g�	�e���C2���A$mO�#�C��@	�*Q��y��l?�ִn�!��Rle�k%ܩ�6�'���,�`J?�W4�;��P�����F� n��I��g�s>�R7�w������`w�[i5�`-Y�c�F$��"�ϣH�|��1_���P�jEC��D5�qXٸ��}ÜH��n�:PU�Fᨕ#��=-j�p�C�4*o��1}����9�ʺ�543[�u��>�����b���P�g�~ ��3�3�zy��H��#�����"@�)��w�_�NS��S%�����^��z�g xJ�V�ݏ�ʄ����C[�dPS�cW�:�G��`W�7#'��@+9^n�@�9.9މ?n/����
����U��d=��[��,��It���}TҝV�"A���G#�ա�V���gD�ʎ�)�=K37sS��,���B��qaF�y�"rf�NR"�uK#�S�M�'��C4E��o��%�
��}̼��v��\�gp�&DC>�u>�g_n�΂��5ߊ8^/˥t����؀�CUx�z0�����9%����1j���]��\���m ��kn3c6T.�]�Ԝ���zt�1w٥��O	@X�d�L�A;��VW+������t�Q���m�40��&�lm���r�9���Б��Iۋ�ue~e��QK�R!3E�k�м�X�x��nf;���b�=xK�k�wbZl�.qs5�����r���}!aj؅Q��H�Ӣ����@���<�kK�x
�u��`�3-.¹��ϣ���G��Ki8u	A�-���Y���U~nw?��a��GB�\�d>dhX�GW�pIt���>�'�䐶�Tc���VB��!��\++u�@#Wnw���H=�ƢN"z�P��z֐���|�o��h�G��6i�ʴ��sf���_.�׊�#@ڄwR�f~y�Ng���^O#yO���Ia����$�q��!r�x�s>��O='��f��ѓk�(4�Ş��j�`;>b��Yk� ��癛d����dnV�����ii�o�o�J�T蟐\�m�:�|�����$���r�N#��K/2�PPa����p�Y�Y��S,�i>j���$�rX��GҌ!�dW�����kZ��DvM��r���.P��?�TYSg]�boas��jګ#^',��'"�X�4*�<ڍ�.z�ݐO+Q��M1X�C��̾6*�x�<�f�Q&+~�	-Hs��q��nZp�W���Y"}���_�b���~=f��&��>�f��O(��%n{r�_�m[�
nE�&4Y.J�nB"�KL+{����{ �ĉy��Y���®o*�ڞ2$�QQ��'�6�ۙu3���y�ș�L)�V����J�s���C���fm��G��2�FR��ޞ���fw�$6 A҂�����c�_y�qD�` ���f�\�ڞ�b*��f�q��E��Npl�	�<a�7�9Q�>�ɐ�\�u���ǥ�39(���O���a/����'�<�,�n�0�BL�"�g��[�/�1�d�B�;&�y�)n!�������1�$lCܱ�9l�-�ϴ�\fF�ƨ��K��P:w����jJ�h�k������0�+����f��ũ �`��9�P�@���Z�߼�葫0W Y����a�&+���$��FKW��BH�ӿ�RV $�M݃��J8L� В�n#�=Tm,QP��[�s��=iշo{dT0d�L�y����N� ��8����NL�r�%��c�u�����#yX�r��8	��T{w=��׌�nq�a��� ��N3�DWN�W�KY�^�:5��F��u�){!������P��ZΖ�s�t��8m��������gk]�""����tQ�P#75��g���^�ޖ̱.9�)��� &��Β]�8�z_08ņ$f
�*^o[��3�M����n��+י�B�#��S�'���,�q�3��@J�O��|���wU��;�)��B� &(��OD����l��m���ve7f�=�WBQ�!A����ep����1�^9�)�=5 ד�C���UX���ȥ�@T�z���4���
�(Wa޼X�4�]�k�D�����T`o\F$��HQ_|�I�?�p��%������d+t�ǘ�fm�/^5Z�"���60Y�5���
�V쏭	G,H��jM�	BNQ���P�����/V����U�1S�pƂ���tF�(Li���24�e9ٶT,���Y٨��x�q���p���v_eR4GHg�?kӂ��}8�1�}\�f8����Uv��!h� ��!���K��;\�!C����AX�+F���o/��{t	�>�W���+]X(;����&|Q�txj���m�MNi;��)�)p��o�I�kD�2��<� �؂��Q�=����(���氖U ���~����jT\���c��Ϡ,(q��Dί��:���_�=�u�/��<�u����#+U���Op���}��ڲ#W_4��ޮ+]w���H�M�g�}��v]�|!�Rd�0lXq���D]�Y��f^���CB(vh�B�g�����"���Nx��	��А�y�];���[��c�9�M�|.����JdX��Xy����槃	�X��g*	,���MA	icaE��@/l�M��Ǒc�!�:�.�9y"a���'��4��ఁ��h���x�:� f��8����ִ��˴`yec���@�؇�'�J#W��+�:�㾦Fr }��)��V<.hU ���ʯ�޻�0�xO:|hi�yy��KQ�*����a���߷ii�Tm!��s0��	PҴ�ʱ��AE���m5#2(B��.�x_�	��<c�W����BY>���.a%F%��%\ 0�|�� ��PS� n��<�w;���I��C��s�8��P9T�]t4�>߫Q^)��#�њ������.��&����<tHqd/�F8g�T���
�l$NY�a3=��������*��I�+�>P'�n_Sp���&���`����D0y���Œ*3�Ί����q��eq���aʟxB�W|^�bs\a^%�u��.��!�c������¬&���&�U�lf��.!c�e��f�&P`��d�����Gv{�VT'����R��џf12�N ZbV��I,uN�����	��(>�Q�=�+C�{r,���j#V���;��x���*��'������ �J�sx��# �S�����=!�QR
����#���$����d�Jr^�X�g�)�Jk�����/W +X:9\���ݲg�c \p�����ƒ�.�6bI�_�d�PFx�Z��x��Y��#n_8V������ɼ�)�l�k��-W�z�^� ������}������R��H�[H���3�/�_���j�<�U�⿒�u~#'��_D�Q�A`���J��iA݉�ϝ<�L@V˨���/]��� m�c������>vhE� 
4�m(�T2�Cj�ސ�x=�2�9<{T">z}N�S�2)����y��p���:�L>��_l�����@:���B���x(��Q	�Z�A��vk���7�F"3���_lN�s�3�:��{+;�%��vςQ6��wdWy
�TmFn!�ev�&��J" c=sz+���]/�}�kN-K'�{��W�{�=�F0���v�D�jٟ�5`t���\M��3���=2Uɠ��X[61 C���Y/�h�$j�寭��J�:��|V���0���dz�ЅJ�Wkh��	�*tR�q�
k^Q�U��$�Ԉ7����N�>Fx�����ȉɣ���ܺ��T������Z\�a.˰��_��e�R��ߤ�C���6\�T������=�Y���/#��|�W�+ϿS0��l|CIc�(���>���O�o�PC_�<ڍ`�1��V�&Za�Y�m�cp���Nt>�˵�MŽ��cq�]��͙F�$��5B�,Q�-��<�	L��'9=Õ�<�o�j�n:�;Θ?[ͅ����?\��0�w��9cG��LTa��P��X��&�3IM1��uZ�hd9�j؛ҨҀ5��*��������xy���j���݂�M�h�����D������C�\G� ����n����0hـ⩅"�&�y��t2�Q�0�Ry�O����}Qm����%�J����ٛb˄	b�b��n*��S (<<�X��J����R���Ґ_X��A}˰b����T.j��`����#܊���b��� ��F�㯩��h�Bܩi�%�ށ�H6�{dR�Jt�Y�U���'Kms�"���n����'4���]wۯz�w� ͚˪�F����#ޞO�ID�� 7�
�?\���a��X)���ֲQ������O��
.�	ʓ��e��uщ�r��!����P:�P����5H�j$9�6(�.�h�~Af���w�)�4w}Amc�^�>��tU�Z�6��]��y/oӯ�[�̑W肧���A����=OK����H�\��_@;P���br����A8�����
{P���V�]jd���VC$m���[ȁ%H[��~"��P�];�ն���Z���\]55R�U0��t��Gx-�R�_��E�qm�o^��*�<��5,CR��K	�=YЙ��F����'ta�q����nB�kx=;h�K�ݙp��CCO08~�G
o���?���"3u@�Y�2�'�T!�oH�MU�����Y�s+.�����&��8,�ՠU/X��+>[��,�5<V��8"���E3���a���b����Ʊ�{��B�������##O���ь�
%!A�N��$~i�|�#��Nw��b��G�����D�{I#�^���k���Ԇ9 *�<P	�iü��:���r*;�eDn�[q�~OO|�6����y6�HrպR�YE���C�{�rI�*�b�NU������Hd̜X6B�@�s������y����	K��C��昻?�U�ʰǛ�Ct}�{w�V2�8�cO�V;_C�}��F��~n��kB��l��
�fp�ra�*h�մC�0����,Gv3�v,����GG��!\đMd Pw����eh�� /!����a��wB����&g?:Zt����j&/|0a��`�����.!wsM��X�揷T�N��GS#P|�_a_�
���n��R�e�y���6V	�X�Q�$�����?�a�h"��t/y�w�$E�1�ˢAĥ���,~�`��>��U��$f��1����~�����܎ʜ��H��*�d`�"F�)s����R�(jYup,���M�����x�pio(��m���{�C�y+iz|F�Q��E������)A)����������CG�8��`D��L��RIw�iy��`�����h���"�Xj"D��M�p��q�*�[|���%�%0Z��`��|�@h@�^}��{Pa6���֊Q�R���G/�Ұ��S�'�J��ܼݲ`]ITj�U��׼h��h��mG�C
�{��I�kL�V}�i0��Q�?]�P���*��XQ�N���`rwdDA����_n������a(*t��{�}K�V#��:NPL�a�%Ze�﨤Es�a��V�6�Fؤ��;X/�2�`3���_�YL�9!qO���z4�M`$]�҈ȏO���"Mdf>��;�����#�G�b.���<��&c�l=��d<��a��>F�]�������� �u���6�������W�Hh/{��z�Ä&�����/9���Ց�gD	���;��,[��P���i����G���;tp{9B����j�<�v��>�/��������Ai�\��Jn�ϐWnM��@��V�Aj1�b���n����[ ����R�m;f��Gѹ��19$k��9`�ɕ�&���h��FvD�F/��{Q�}D���DӨS�f83%�)� �3��q�O+�{5���BQ�g�_b�B%����(���(�Vt<K�p��)*�B���Q�-FS:ކD�ip߈�l�P��@�G9!�mʏ=|'9�oy�9ǆ�e�D��'�U���p.�? 9�Q���c���\���W0�;�@T�}C���7	U�艄
��ү�L�9k��[̓~5y��آ_T�d�+�KHH���	Zk�oJ�[H�bդ���-7���/�Z��Nid�Rn�K#7_��w��A�%�+fL!X�Byۿ�p���0Gk����|���c�MW��{
�m�Pc��H�lH L��9F$��X��HG�	��af7ny�q=��3u�18�O���q`��!�a��=Q.nHq �Rq��B�%S���9)�M�x�~����DD���y$�&�D�i�����FXK����~�߾�G4Oe�;��p]��J��}�;ǡy�� ����h���C���
@N�x>&c���d:U)\�P�m=�@�S u_
k��7��%����.�h�|h
��ut��ﶄ{EPy9یS(X�b��y���ʇh��%�|��读��9�z����b.��:����E1G���[�~!Nɚ+:�g�7�C�F�@'�4�'���Ρ��ؚ�b������B��+09�cG�Fr����g���ͻ�D�%��r��������ʂ,�vL�>��J��f	z���(����*�m
v6��O���;ڝ��$�wD�ܚE���_��+�����G����fh����n�@m<x$��0D���#H��i�y�YV=Y�?~:[�L��=7�5��PGt�3���V��T����~u�bيB���%dϿ�d\�K�[b�
�Ȫ$���{���-��4A���9O�h3�ZU���a��z���w�<��3��r �2����f���ȭ�Ғ*�f���{(n�<n����=���`�ր��S�B���� e����c�6%8�a6�(1�0�ܶ:�OX!7o����n+@L����������r?�"S��ؙt3�|�k	��T>V��#�Ŧ�5缒� +��?`��_Y��)����0A�c-r*7K��[{��@�?,�Wr�U��V4�!�p���ۥ���W∼"�e�����z.r�rإ5���pi	�e��p�'�&�4��ۡ_0��a~2���<h&��hfTa��1��[�#��R+���(�_��
M~J���b!��]�d�(�&��TCS��퉙����C93g��B�N᫿���C�쁊`Go,�e�C��v{ڲ 6U(��i6l#�e���],�����}d�����t�gaM&}�������;x-��y��]��c=�H���,c�FD��[3=81x�^�����9y=#K�_E����l����a�,	��V�)g�s�[��I�H��У�gd1[q����ٍ���G�}�F(�1��m,U Y��li<39ȔK�u�7z_���?��t�Xn�!��o��R��[�G��1��G���>���S���������I��%,Kj\�#o]3qXUn��J���������o$��H�M�=ގK9U�a5>U��w�D"����9��T�$�iI�D�B"�>��9�.ۢ�mE$��7��~��]�9�}�[�(�z#��A���]S�B^��#���^��9;W��Kd�d0gN��.v���z)��ş��u��yJ
�9��$J�23���MD3�>�8'�tc���ڈ��,ɘL�~u���F)V���� ���.d�� �o٧?�������\��c,����ֱ��ˉ�lO�;�~�C}!���W�ݺ�8L.�1#�λ�6��x1�M�vB{$��5jT��Up����(K����i���I716Ұ� �PW�3�O`ފ�([ɱ��h5�yX��	���[c	�N�$n�.~�NY%�=��V���ʶ��ڊ�
vZ���#��3��n^!��q�٬��K�x�"�2<��z3]�<�*��|��r��ٜ�i�猻�MM2�����Bq�,3�T�1\4�)|�G�<.'�5yRE[Y�Յ�q�d�+�T�C��Rkf�p{��~5�U��ܗӽ"�w4DB��ժ �Lm�B!i��#�l6<&TݝO�J7�1�"�-�qHU�re�ׇ&�((�	DW�LXS�2@��Q'`M�C��YTIJ����mV��g�0Th�b�������^���[n���e�~U�WI	 ���J��:}����[�?��A���/� �Z_D�o�j�xL -_�T��ѐ���C��VP��
� �>RM)`��;
6�HRsp�zX��$�j��'���ܟ
���fӏ���-��;0�a���m����ƣ۶�kZ���#2%@9��zx㺰8���{�F����]M��J��띨�̓�b�S����[h���F�m�@H1���bRTX.ݣ����bP�;o���~
k�J�s��C{#H�2��oJ����1J�숻�JR$�n������ս�\��F���U�]|��\�� ����&g�,^��a���ƨ�朇ܥv��Ʃe$ 2uҠ�uC�w�8���%d�/����m�]��ޖsa��O��w/	��W-�⡺��^��觶�L�|��'"�+z���$��q�v�|�W��$�G�A�
�GH�Y
�ip�\%E�Q���sXG�[�xw���<OGl�Jx|�B��!+�)cO"HW�����X�cA�3��V����[���vԙս�*��������T	`&E~1<hŧ_�����F}�YI�.\�a>�?"���$�aX\�ų�l[.��*��##����{�6<���+]�a���tl��)M��Ә�7�3��jm/"��PC�d}�a���T*�{��o��sA��=���#!�k���w�i����b�	6ڟ���@�D��U�͒_���6f&����S)T��L�駴ٔx�#�)���]gy���U�n�<������u;��_�����/v�؇z��:j��%a�:Eo��]��6��_�Y��g=`���B�Р���}wc�<�/^v����l*���Z�W����T�n��fG�+�{���r���q0�$�	�\rj��nDn�����Q���@�&�Wp� O�����H��J�U�Av��T��>P�Ľǚ��NϝX��_zj@@��J$����;A��H��<¬�+� �-��9����=��0tZ���t�|��M�ݝN�T3J�!�/�S:о��@�"x��$�f)�0L���EC�8��k;6�Q�O��2�v�mq@_W�gNf����}J�I&v:��t�,$���\Z�u'<��V��'h눷�o�Ǧh	��!߈�~�y�;�d�JT^`��c�#4nRMC.47d�>���iM^��L��(V6>��i�;�������u���T�)�C���sͱ��� ����QC�����}jI�B���tN�{r�Rc_���.m	rD;��W���ܲ�-����L��Z~'�|c�~l��bIėK?�M��v���Ծ���H�Ƚ�M׼����&䌀����v+�Y��t_w
̀@ɠ����>u�%�f��m���d�����Dn(�<�Ns=���d(=�
z
|���i�OD����F��^��!?�|M�V�|��3�4�0�D���O�uj�o�`*�q�m��֢��R�pI�Ax��5�"��6�@%�s��uRW�!�zo*�;R��F3���Y-V׾����ݹ��֚��*wAauN)�O��[�J���}�/�Ψ�_W_� 7E���J��ԴO�,`bA�C�ksR�YI֯Ї��C��mށeJ~�.eJ��pJT�lk���=�W�����zX�z��|���S�)��kti�����GD嶐�����J�Ώ��O޿�8�G�m`�7�gX';�R�&���IJ���t�z��{�� a�4ꡤ�W_�s���[NJ�Ed��}Pֿ��Y,�G�l����[mx~�F۞���� j�w�����qU�Jt���+��gu�~��d>��(\�����A�@�c�#����(��б}J�e[j1���`cU��u�fw�#�]GV�`K�����+p��9OG�|��`����w\ܥ�B&hGRnk�ۆ�R6� j�]�ph��(�J��*�n�`��hP=�(Ӈ���&%��^����[�=AW��)��ʱ4��R�������ס�������n+nA��B�bWR7���ݖо��x�ۂ܊^]%��DA��+蔴��lȚC����B�!�NW~T�p>a�N����!�@}�7������%��g��/-FǊ�d,����� gR�.�.<�v�}/c��D�%\Oď{5�4��(���Y�Jٌb��!~�g�xU�+�5�(4�ψ!��k(�Q�&M���f�^f8�G*�I���V���dEN�#�b��#�s�}�uS숚��V�}D����?0�pn��̪�D1�$r�j$��K�T�����{��	�t���8$������|<����_|���M��/�W�M��B~ ��[g��XXtT*]����,��h�j�I�u��ߥ��@*�K�����#�z��U��x�p��Z��#�kY����F�bP{�7��a��&����4N`�t�ff��v�N�d�.�c��}�&8u�N�>}�����SCK��LM�X��N�����"_���	]�<?�N���&,و��v�����!j �P�����WB}O�'=�ΈO�V��˜�;�:51Y�����&o�S�E,G�z��y&Iּ��p�@ݻ
0�?�E��-�S�K??iT^Z�Y�@�?)�Ut`�W�PƖ����� R��m0�g�!�欛�nn��9W�7�ϼ=-���!& �/ 峤��U�lS?�s����`4�R/ǲ�~C�[ }�M��8���e�\�Yj_�^r3����j�G�?����U�8/$c�r�μ�Rط�R�b�[%���jk�3ꤸ<������V�����b�ִD�v�����d7���v>D7AcVC@f���^ �VI$x��G������T*:�ϣ9��l���r}f޷�g�1�#o�޿�:�" h���a3q��
�@/j�,M+n\��������>iQs(Q7����6.E%���(�f
6Nd�Ҵ��銚�W@�h�E��@~	�
����_(~{�Ѳ��n�d��L�˰j�����I�Y��2��Z���#�e�?��S���U��J��Q S&��cǹ���Q�2�s��r73p��l/�!8���H��R�{pS�02����U��NG��jI V����� �vX1��64��ai���S��|V�9w�lR��z���7|��!Y�̋����[X���.ޓ����2Vq���ȹ����:s.J��ڊ�-�{V�����]�2t��&T}���S�䤈��꧀�V���!��r:��`&ܒR���ԃey�l t��ĘV�M���EZ���ƻ�u�XT<'�\rZA4�� ��#V%��si :|����*��&Tq��я���'��tOl���7.pdV�o 8����c=��O}L�_�8uHQ�0��Hh� 3I��x�� "ݗ��z���a7
=s�nb��M�}ԙ�h��kf��40`V`MeDD,^@&���G��o�N{�<Ю�3T�%��v��
���p�P�� �Y�9�C���g��VM��g�тm��]��Rz�l�5�d��ۗ����t��Ï���� ��S�n	��Ho����֥L�_kÝ��\,y"#EWx�� ����4.���f�'�����lu�W��u�t4L�A��F`kG;ko8�3;=��.��Vpe�2;���x���P��Ǿ��,�����b���҉f��:��֍��}B<��B���z�B�+���8�g��]: �*�~9ɽ�\��3���k|���<3qo�QH*�����t^�`������E䂌/qn���Wx{��q�f]�����*��x`tV/w���A�K�?<F�1p��>l6vJ@�@IhGɢx^� &z����8%{%-���Cy�֝�d/��~�hr|��ֵ^����A�>>�g���&�w^�&|�:f}���fM0�n�q�	��|��*�����e+�����v��N�q�D�A����<v���Y���ݮ��e��Y+,�rC�0B.�:��G��"L���3��3�o���s���U�@m�m1��P����C��R׆{"���n�z�����m�E�D�+/�A6���B����=x�i`��W����	�k�J�B�\���l��%oo�݂�ϛ.�� ���b]Z8�
ʀ.Y�֦R���yJ����4�X��nuQD2�Y���[��j�cL�]HN'�0���H�s�����3�:p��	���v]�xj������%	�\N+&����L*7�&CQ)�F��~���n�E�ĎY,b��H����a?-*��^����(�yz���*��&�y��8�]qf\S�fJ�3�o����B�H;�"��F�;Y�R>�h��^��lH�=TLy�|ɔ��	����6P5+��[kl��� �u�Uݛa�t&Q9|	u?�䭞(�<G�9B�m�:�~����Zn�
v��s������w����[s��Ί����Z^���#@)��t���j4}�Sx�}K$���v�;��?�.�fO�w�,C#��,��T<���r��I�3ڊ 
�����ߏd�����)�����[�:�i�:���Ày��+X(���I/�pl��9Zq
FY��ֈg����L�}����UN���%�Kb#���QR��S`e���jXM���p�w���M��e�ѐ"�#+M]	� K��
B��_��_�<cd8�#�@`?�԰w����h�n��Q�v����x�ώ8)��0R�lz�L.}�������¿�<�������\釙E��"/������x�� e�e]]�k�������o>�θr�n�c�T�\1�)f�k/�Mg�m��U5
�/�,gf�/�b�͔uf�c6Yȁǟ������@��	�z����2���K[�o�pĂt��[���tU��� ���WeJҮ4�و@��C�D��X⡷��hB���˹��-�i���ܼ�~��\`^�=q���c�z\��D����d�vLYd)���Iz#�߭��j�̼P���^���}|��{_�����ܓ�F�+#��`�޸�[�� ��$sC���o��_pD/�;E�ت�,�}"� �Ig-pM����I�@�����|��d���4�����D��r�,2�������7���g�N�t�:͎^M8ټ�0�ۑ�=�e]9�L��Rv�*h;��
q����*٣���ɇ:Dg�iI(��p�΍�;8䡿��i"���U$ ��'?�o��pT�a���1�Y⪺�	����X �#�Pvظ��3�s��{�^&�5�֟-�0�V"�9�i�b&�V} �Q�r*纻���ˊ;�҈}��?�ߨ�IJ@TEcqs�]��׫�f��s+S���ߦ�_���]�('�s0L�H���|
��-���^�&ҩ*ޗ6�=����	������yj{�E盓Y��I�m/�oi	�K��
���nL��Aq�h~�a�#��dd��o_��T��0��)ĎF���c�T�o�H-��%ec^ ���4BV���9`�Ū��Nξ���}��d�{�g����8�a�ޤZ3v�>������(�c�(�c|_�2�\pD���E�|�h�ZG	����I��y���.�m^�5��A�����t�h<i�f!m`�Q!���K���r�r�~5��Pף��*��&(ֵ&���r�-��� ���?؅����(y]��h��wxD���o\r|d�ORW&�>\:��ЭZ�_�vA��}iK#�n
���A�O./�͇�jЌ�cu�!ڎ�{��+X���d[P �7���Eq�DR�nL��t�����#7{j�w[Ǘ��14�!5f>7Ν�jh�gKthz1@��
�� ��\5Q";5�����e�{����w!����i�Ν�e��J����.��N�mP�&chؔ�T�#CN��N`�
�RȢ)����=��:�)��($��_�e�K�vX�I�~)VA1H~������q��\��1P:��H�$�F½��ѻ�U iL�C����s)+�}��o�Y�WUَz�-1�NX�N���	ھ_�0s"��.Z�x������sa���?R�0��
��BK}�ԗ�]���,�ҙ�����]=C�,ß�jv*�%��V������}��䇼-�7��AD�p}y
Wp����o����o�����>��F[�K)�pD������è�����o���ۂr+�[�v~��a���ғ@_�`�n�m��Xr}�.�$3U/O[\����3-dZ����^��pz}��HԥxyE�=��df����Yș/��fL��ﯨ�)џ�C5*�Pmϻ�bRdx �)��`ͷ�ǌ�k�~%�~�$N㸂*c����(�!�(�Q�h,k?'�	�U{��I�rtj�[n>�vS}�mW�u�+��)�X6HB{�N�U|���!��|�H,~I�}�aۘƼk��{e���G\��G�4��p�"���f5RX���!x�چ�\a� ���ܓ��\�#��5��)nfQUG��(�ϛ��)�(_��d'W�x�RR�6����Jx��y+|%
|B�m�W��X�3�F^�`hI�:k�$�=�I^������.M��kÚ�ąٓ�"�
��=̅��=��c�ӂQ;O@��/7��W� lu�}�[m�ġV��g���0�����&�9r�s שk���`�}��3M@�KU�aޏ�P5\�o�vH��	X��u��E����-�&��_<���ObC���+�$掼ʺ$&�pj��_�m��>��a�z"����D�&��Eł��>����/Q��Џ �����ΡJ���lh�H�b���ܷª�JS�6�B������9��n;����ZI�
vN�;����PpǇ��O�}zA� >�U�뽣��Ny�?M����-��G�ž�Is������
r�t��1�*��p�Ӕ �x8-��gF^���''�M�[^�o4����N�-q�}��2��>�<��t�J.imߡ�Un��nεQx������Yg�*�M��B�(W�^���-��ٖ���qS�O�Ayi"��d}�j��M[��L!9��%_���i
�����fMsQ�̕B?�+���������ѯ�C��*�=4B=�t6��s9��4cr�S��.�r��Ƹ�vX5��ȡ-�崊��=c���W��C�DE��Sm�B��~ ;DWg��v�x��2>`��yZY��Ui�-WSQfQ/4ޯf������F�{�XMRpxء���������ƥ���q�A�Mt�]���T��v/��pnG�j��F�Y��>V4� &�j2�FU�����b��m��r&�¡�?δ��']0l�� �zO�X`Vձ��%.�����q��*�(d�Hh`�t��0��-f4y�ͽ':�}>oO�*^T���;�V��=���x�'~�vOS�(�痝��؄�#��-�l��b���;^�W�nQJ��] ��}M+�_��0��� �薯��M�b+B6�u1��M�i�Z�q4T�&�IVZ�V߸���N����;��~��>xSY%�[��owTr��ՇnSb�N1s�ޡ��6��NF�b�y<��A v1�} 'É�����zZ�]2~�z�k��O�V��=Ǝ�Y��/��}���-cCQ	����!mY���q	G�Id��ݰ����ݛK���hB;V5/����y�*�o1��4[����x���F��6o̧��[���'T4[2��W-��*���ą���m�%m�@xG��PD�a�!X��\�R}ӿ2�����>����4��-�:k��	z�X�>6��L�Aڌ�!Y��π�}@�E*�c�@c����(r�<����uz٨�!{JSn�-�x�hv.���Ѧ�?���%ġm�ٹ��-����M��IH�ܛ]EB���6&ֶ�!��!ٛB��6��oj�7��G0�(W {
X2�|pW�*V��Ͽ�t�T�~�\���p���4��M�Y�?��7��`����j4�[���#ftq�x�M{{��.��������Ni��ݲ���|���
�o���1GJ�,!T��ڳ��]tJ��������-n�����OچO��M�/DкQ�ۨ����52"��B��>!}Oc|шř�<�$��h8���[���IϠ)x9�w��!-��ߛ���������<����r&��kB��z*G������l��˔�����Z&;]Џ���|��,�|�LZ����.�q�T2c��(��_z�bX��Xr��������ٚr���\�Ǯ�I�[�/�W/����!!���;g�J�G1���Op�o]�Ug�	�HhFW�ɛV�֛�����C�k��D����<[�x1��#��sM+k��\���%�'��(h���?���p޽w��=�^-b_�<'���aI;d�z���G=\5�p-����4�������8����I�������GJ���ݫ�eg����8P}$Ӈqu�}��o)��`�˲m�<�<��p%���E����2Cej ����!^�{�1Jk����ݫ�5lxޑ�xM�q'*���6o�����?�U)J�5�$���..��lAw9���c�F��~�� :�Dٌ)�/��g���ARu�����F*����y�m�W���n)�)y<pT��:U�
bF�؃ه�էU�|���.�k8դU4���*�M�&-Ԯ���	�t5�N�D߮&�SǗ��O��w��W�l��7�lܷ_�)� 	�k��e�{����=����<�x�_ i�ݥ�7���'� ��@*)X��ݽH�u`�Ǖ-���
�[����_TM;�#v��脏u�	c�:U����*��\$l�d�J�~�#��f5��|[2��������,�`���a���k�ų8����Ek^C��"��wi��<Z*"�/���,�O����|�z�nm�������f�)�g7�5�>��01�Xi�ihWNL�U��9R��o��ז4�x���f�84���>7M�>��'��s����;�g�*�o8HA��M`�8���_Rp�0^��W�z�6mzK��H_�l�k��?���c��qv)���t���p{��آ����&d���]t��ـ��ʐ{���S�]���<JK.-%W�Wa���)��F�a���y�9rzU��3����W9�ҋ.�������s�#p���&�+�)�<�wٍ�?1����@. ����
�dӧ���j;��)�V�����=��C�dc����kC��V�Ʌƿ�7��-X�J�o�u.���h���ҡ��Vg���=Q�wfH@��.ecXΖ뽵?��[�Ȓ�ΧN��� }�8�v��y���6���P�h��� -Q�T߹<<�8%����R�wyS1s�g�g�l��%H	�/}KVs$�'$ׇ.�Pt`�!1d)/�:�� �`8� � ��waf@��A��'v�5F�m� ��h�Dgz)�.��#�\����o�t1uik�j=�|}�-��/i+9�����_�U#Vas=$LK�Q������b��!��hN�� Z��PV�뿵?=����= Fo�J(~բ���9���g)���{�0д������뚻�2�ōS	��ЏG�2�D)��y�oh�{����-����5�j1ȁ�wg��vqZ�]���;�?�� U=R����eN�r&hj�^ͩ�$��Sa�9x'���~���:?L{7�<�h<��i�ys�~qf��G@}vA�"h����稜���^L��2�I����A@.��!�P��=�#�$~�h1_KX�;�(��C]m��a��(����l�����|4�L5d��?`w*��)i-m�<��ŋ��������Io�Gz�jQt���'OMbԄ�����#������a����KBS������́�K������+^����G�#l��醂v5XP�����̭RuSc�[�� �vg��Q�ϸ7���]x�[)�n5
+v�"�� ��j�ϟ�ʉ�dE����9k��̅�4t����f����~��T�s'u 4ž��~�cc�ǝ����Y�~�9l�Tl��r�J�HMd�>>���=���M�>C��АX5)D���֚��"����ѩ2��Ԃ}�C8�^ˑ�v	�(�O���5���&G�1lT���t����z`z���a��HSV�)M	�'7��f��()v*��1���PjׇQ����
L����>�5�^l�;���1�NUЫF`���&���!����c��$��1'���l�+�SM\���M��/�[�G�[���+�[�Զ"�)z>_��X\��I�_�ܐ��J@�\o�Wس�$�uD^!�î�|gV�j�Q�<�Y ��V,�x���IA�Ȑ�b��� pd��t��_�59N���-����g����5�ݦ����7��3�.?�� �B�qխkFIFl}^�S.���5́׮6
I4�Pw	+/5�QjR�)
���x�,2��>t
�����2}��Jǻ����``�9D��~�����4�&��]�P	U_6���%Kg$�iҙ��ɬv-g����ˣE9v{����}�ti}�r뺺$=�����l���M��4�y�	'ɜi�h߲DGҭ�$���IF��]dY2:z���x�x��Z�*#Qp([�"�q�LK�c����:F�#x=<�)�1ζ���l�L�?2��.V�쁮z�ٖ�"Un4�wC�V�t����5LL���P2�y�"�v�xSEާ2��.�x�[��_2i<z���G���4��I^G��|���3��c0�ཞ��P^Z�+8^����]�[gϙ9as5P{eP�:
�_�Z���]-��fstR�i��rN 5F��(�0?��J�ӑ���=U=��'�됚���;4�\ �r1塗�/~�]ubW�{�(���ZQ�7�����g�A�dik��y���Ap%`�B�aN���S��m"1���r��M���|����b|����/��כ�Y<9J��I��M�R���~�Uj�n��ݵhE[���O�?�^]5ۖ�:��&d��Rr�$"N��-���_2lӭdK�5g��Q�]d�l9<���֦�
����z�+�ݣ���z�픴j&7$ށ0�845e�S�`7��宯�\�kȔv����h�=W�PFy�I��S[v������T5]�J�Ma��N���~�p�(�;Q9��$�B�����F
����ne��wS"���9_EbFY���{�����r'�\c�
5��[8�R1�B'��*ծ�(��j�>�?Z̹�~	�j�68%�sh�IM(_a��U;zj
`R>�:�߬�8j���z���$Kv
�t��w�s5%B`Q�-�n*��(BG˳I��2��J��� ���{]�nOI�^����0�_,���Op�*-#X/�3K��{Cǭ:�"Y���#������#:�����]�L2�Ow��5Ћ��\)9�L��a��`�ٞ�V��mæ��N�"�<P���T���V�]2��JJgp�2�^��@�'�Z~~M�J#���j	��qܾ]{��qw�&�|.��i�}=����H��E�v�$.{^#����x������
���by�����i����<�PRϑ�$�C�� ��y����**Yp�:�Hj����St0�b�f��	H��W~�m��c�DN�eK���W��= cw���eK(d�t.�`����|�!�a�i���)6�}�k����8���RZ{֍i[�+Y�t"~
�2����fV���Yd�)D�.�ߨ�y���ԕ�x+�v<��JD�ֵJ�G�d|� �[8���Q7�=H�l�W#R���%��>�D��4P�I���]v"��}�"Wp��~�N�̘r<F�vob��*g>���g��W�]�UZ���Lh��MX��I���������X�š���'�4��@Ir��ֳ}*���=���*��e�ϜPB|2<;\���n"�S�
��_W�|+���^�E
$��s�}�-:�	m[�֠"Gy��py�54�9t*LS]N�e
F���, �b�q�t�A V�*���|g��!��Sl�p�B������M��1�� �e�3�`E�����u�o&�͂�@��@����/#*nn�G����)��gv~Y&��v+�%o�q
B����+*Kv��]�v�c��Y�������)���txW�\o�n�r_��񤈐�"�9�}���SNP�������1SA y�m q��.�V��/�>N���h�M�~�5�K�{���;5֣��8 �/�-R���/���n��ٱu���תP���fR��5	����yr�M�a:�Kנ�����~��n�Ct/'%�\K�z�Y5�H(�,N�\�uK%Ik�s��P�;ś��p.��>��d�4�� [3�w�kmȑ�~�l=���TI��2L�1J�%s>�Pͺɔza�����y�?IѶm��k$�>�ո{q�a��F�M�-܃�ڲІ����������Iu<XaW!�J��W��H�'�b��kz�Z;�bT�b���O�(�@q~�T.ŀs�>��a���ڮ�+�9�ŕ�j�r�_�)<uߡv];�*R;�"D��w̪�7L��Ƙ����������⸌����z�E�T�a 8�2A٘���\u��e:6o�5sK�6a����y,�ՔZ�Q�t]�����o���J��$�*��v4.����%�_�'~ߵ/Q��ea���$��hsF%hg�0�F�#S����dz%TyRC�`E��������r;��Ӏxz����;�M�,a���Y���ÈK�
��"�X�k�ٽA���Q��t��+�'u	H���=�v�؜�!b�Ae�;��U�X|SHw.���wC���ȩ� �5Vs�(�����=;��Du^1�R�oG���\�Zö�_��;�!�i��	!œQeB���K���t��P��4wKT�LB���vT!�D+Y���g����%���(�o��k���?�GY^揃kx�O�����`�cĦ��\����$�R�37�
����XB!	f�7��x�2�;����hS�YD�|�!�����_�-��(���pJ��6�ͨ�ig}O��>�~�ys��+�sY2��-�yad(�m�'[�Q&h���2 ��j�j�!���Q*e!�x*k�t5v���O��gj�ի�<�ϣ�ֈ'���z�*��#	M�ӌٮ�����K�gRj�+�/`G.��}�(��Ҡ��:/a_��i;M#뢖uW���c��҂��J��~���nY`	ahV�"�"�b��(GLs꠆[xj������_��I�%ߗ��5p�\�o���b
�1MԊ#����9䍏C�����A����6��n�gW�N5$=K̈�5v$��S�� g{Q)|�l�#�9]�?��y���Fv��/�.�"���'��׾�)s�PF�#�g�$!��J%Ko��K�v�@�1�Lk��q��H01��f8f�j��Wc��*!��u(��c��ǖ���7�i���*�����;�Y�~r�)󆹼3�{��:�"?�qc�	���U�>s��d��[�Q�G�s6������xi�!ϛ��kX��O�~Z�;.�ty��e�P],#�3�Y[�w}��J]���pIO�����番^�gKV�RU�����obO��Es1�X�V��DH#�iV9���_d�+	@�'O��-
$5X�VA'��*�<��X�(P�w!��|m$�c�@�4���� �8��O#kK��Ns�����SKe��?X8X�����I�k$�(��TS�)�N*f,?�Υ�m�s+(���O�d;��%�A��@��H3�2�{E�8�-�����{��@������Inm���B}��0���O�(nP0�yudrIHv;�������ǒ�dXS.�����0G9�u��ϣ��'����~q�VZG��¼�v� I�C�Ў�!�zוdXmw�C�P.M��g��w�a��&7(��n�T���w�P%�
����a>kTL1g��#(���,o��G# ,nwי�����j�gKݭma���@��I�cR���;v�t�mP�{h�Jy�5�ej.^ɐ��X_n�C~��Q[Cskl9�Z�KXT_};?yjx��cUA��$�f2���;�o)������w#u#JR�@eh�I4s��t��W��/Kp��?/��س��k�fJHg��Ub�꿠�Ŝ��(/e���ͺ]S������-G��DAm<�����<���m���� ��}� ����(�1p'��n��7���"x��w�`�l|�ڢ�n⼃�R��7���?�U����k3�a-�i�����N_R��P��������G<EP��9���e>���#Y��V�7�Y��8�����B��������*q�� �����b	�ݼ��mI^���lk��N4�e���8QR�5�Wζ��f�aʎ���O�0���x�!�8�6d2��v���.7w�Y�%��J������m7_�M{�%���a�R�1ѹÐ�e~<X�W$+�{�O��$�1h�Nֻx䌚{\O �P# zˉ�~tj�,]�~�G�(����T(.���6��[#�j��/�;�����%Zt�Jb�V���FfA-w	X�`�|J^b>�)�/8x�\��JA�1(fM�-��.-�V�x��/�Jp��1�M�s�wz|)+��ً�^IdD��E�B�w��#���6u��:���%3*hL__:�R�8̀��V��]{��b������+, �d��L��^��n��'�́Z6��l|>@�1h
3� �D�z���� �k�3�o]GtV��`�ޤ�>��&K��v�v��T�R��|��9k&��V�m�n���q��^�/���xUZ�;�˛ �!����_Y�4za8�U���Ǎ��h�x �%����>6H�]�h�����
eeB�-y��B|�X[�2�l����n��.�*X�q�4����r�00vK��̦2QG�Z�2e��rٰ\]sJ���I@i�f�O�����r1��L��=��x���k��v�P��ץ���`o��elV�z��HۙX�j����[|����8��E0G��G�cj�%�����C�Jh9�§�f6Lo�J�'10�"A߱����ō��%����ǯo94���P'��XS�d���k�CN�Мc��8 =ޙ l����n/��#i�q����V���d��2y��t�M@k�����:!���Q<�c�6�mM��kx��y�C���kx�$���!�J5T�W�c��/�����*��T�q�ǓN�8n����.�IOo/$^#E�q����I��_��<������<�s�԰��~pP��ՉU$e�����V,���ɺ�-m�ة�wIRܽ8�b���a���|�e��r���u�9(�x�,��1���õ:�b�N�ư}ʠ�D�ͭ�t��m�k1Vn9�X���C�S;D��t���G �WI^�@\�c��s�_`�Ƣ�!�2Sъ�Xik�f�b�pke������@�nK�?��W��ض��n2�['���g;i��[B�	&0�Oj�D�$b^h��0~����RYcX�Ks��\�������n]l6��o-d���1����3k�1�nZ���-��Y�+�Fl� �x��U��d��ތ��E�r�{�΁�]u�㘞S��30���xX2.�~�5�-GB�C�%�U!�)�Lgɦ���,0�'
@G ���3qL2����90�2�R�����5[8��O͌�e�E����4ǥ��qn&�<�&��fF�Sz/�o�s~R[�:![�ʍe���!�ˢ��F�״�@<T��~����1�����j;4iY��됼jm�i�{�����4����}� ��s�T/|z�(�K�1��Ӓ�
�9�T�ء�J]���A�A�%�r�F��|'�ǹW����Ɠ&�	���d����>���TZ��!t[��� za������02ںy���EX���M��V��NMa<�*����}k�O�s0&r5M����i�ai~r
�}����D+��N�F��Dba���lE��%VCB"�^vR�փ�ѓ�:���t4
��Ȃ�2]�O����9#;�	&��4R��Uۗ"k���ՊhZ���~Nk:D���ج}'ϕ��"ݸ�WWcA��;�j��.C;06�Hݘ��e�M�����*q��� ���Ũ�-)��Ƌ=�(��>�qҥ�<�a̾08ڢ��Wt�[��|v\X�AwK�~��WΏ7�И�
'jf����K��Zn=-y��V��I�ZX58��a�ͽ�"��2WZG�܄-��E��//av�A�p�
SY�	�h���U7��H�C�ExY��x(�չ�5~�Zf�eJ�~
Y|S1Zp}k�����,�z�Z���m,!~����ʩ�c'�bhC!��A?\@_`��m��Nմ!�j䧴�e0,�U>��ќVz���Ӌ�5Xv5�@h�N�����Eƺ>��j�X��M��֚���euѣaQ�\j����_ٟ����	^Q����0�Dt�s"�KLx�֫��~3��>�1��H�9�r��ϙ%�5�N��V���/)3R�E���!1�d���X� *��z�~M�"���tt��w<8�c�W��=�2�w�$���>�+=Bu~ߙ[��4Q\o^b˒�V�68�`恇��f�Ŗ�M�:�fx�گf��N�l%y�Q]q�'��W����Һ�4�>��A�DwX�/~fr �D"
�b���JjU�q��*v�Y5��@	C����y�ey?���^D�}0f(��6{`�iϊ�u3���Y!��@�E��{��#ed;S����'�<��.��=k�B�]wKr�ɓ*�+0���g�#��v�G�?Y2kݙh���B����!���l�8�-zZ����j*�U�ci��з��
�hM� W���Z��.��{���x�	�W����J�1�X��=3S�A62���`�LS��C6M`g���,p�Eɇ��� \���<�_�
�X ��`���m�B~لE�ח�Dg�	�C����|�G؃���|ycN�&S��;�Up���:�:�l۰�>�®%�ݜS8 ��k\�!u�(�{���%8v7�sheK!���$��t�a��ܺViX�z�ˬ)�CN�Ʃ5�A�R%��:T��� �Ç�5x3 bőr�u���	H����i�����gE�U,]�j�+^�vD�&�Ń}p�J�l��!�S�%]
�:�l~��6�J���/
+���Oe8"�4(�>���-S��bKQt��b�$VGV��qj�����\�߭��$����5@v���s�.��د2g�Uh�!^�i��bC]�/s>�-��kM�T��o�A�_P}mL^hV�{��,�M�l�lxX_�OۛJʵ��*�w�0s�����\���'.����Qo����ⶋ���7 �6�9tAě�҄.]ZY�2�v���0�݀K4��f�(q�-4��� V�����A���m�� _� S��a��m��r���_�l"�&��T|�=��,��i�i�_�&��h�мQr�c�v�[.�1K��^C5�t�¿��M�V\�2��_�o���vMi��Zz\0�AU�|nu�@�Z���dV�+�d=�%�6�! ��c�Y�G���,�K�8�����R7� �aKL,.�G�{��V��$Y��u�	��d�K��ێ�C9�<Z����W�=�A��en"-�(&�2 ��ɷ�{{τ���kX�g4#�RE"�o3Cg)����"7 ��,�t��<���b��®���ƃ�"���@��`v�	J�CS���YE���:��G�Ȣ��[�4�|�7>�G0���pv��:��n��
�%���I���Bj�twU� uq��$N�x�3ڹ���ݫɲw|�ҭu���n�3����6��u�`��Q=���%���|BAɛq؛�1�'��Y�@#Ra��:� ����c��$3�� B.�}�|�-iXwŞz㭛/lm����6?S�A��?N"���&��bZ�UM0��}�l*(_��f��;0�ggGs�[�Mh |���$,��g(�e�k�)!���rt��WA�(GU��;�EM�_����L�^�P���v�T&L||ng��s�p�A*���SIbo[�Н��;D_K�A"��s�����%��� ��s8��f+�.�j�]C?^n�U<�>_�M��ۣ��=y	~�@� �������MU��1��� ��0�����Ϙ�_)BG�����b*�v��U�f"���# �]��-�'��:/Q�qo����-#�dv̹�'��?����B�mlǢ ��
�)�[ؗ�M2�J���Z����满����߁5|e�#��qO8��8�)w���r�N�����Ư�#�7jC�$��5"2�2o����.mB� �]���a��2�9��20�}�(��<f�܋0g�껃�k��R6�k����bT�#i�:�K8zM���eL�u�0]�U���B�d>oc�v6�:-$O�����f�3�u@_�����͖y�W ��������J�FH��-����A�7y!��5J�A�i__>�sX��K�A8�� |L8.�Z����ʒ��?���4ym{f�Uŝ6/��0Q�0�H%������M&q��	7���'{�w�\~�_`?丅�J��9�XD�7{i� �֚�ȳ�_w^ U��S)��Ɇ��`C�F����*�S��`ߒ��b����9��2�iwš ]�dǭ�>]J�^2�~#�����D
�"sS�sN��q]��)��,��>�.:��ՙ��7@�^�W�`�Ҝ��Ij!="�$�)'Z���ɲ�1#�T����8�)��I°���_<f�7P��A�u��_:{
[���"�kdS��{\�)�3 �pFX���:(��L��$�Y<{�$��;�Wx�j���"�)%:s��G���ք������rh�J���>�H�3�yO7Ʀ&667l�$���yX�5�%	�:�Ţa� ��ū����Z�����P�����v�K1�X�PR��͸�|w�j.��b���3L�4ū��a��H�|��HH'����=(f��B��d��V�/ˮ������~!Ś��[�t?Z�kg��%���U� �A/�)mB���E;�>�SKTPD՟Pf4v�wF9
��yߓ?�	ðp�a��Z"�I�W��^E�痾Ya������W�-�	.�+hՈ١���蚸'Fv��6e�|���J��sZso(�;��b�W� �\]�,cl�24��FY@P��]�q�<+_	�%wV�l����^P�Z�/\���#���`J5/�
2v�A+�d�Ұ�R�Hb=Wn���
1�mB��2�T�fTt �uZ�j6���ZYU�P�d���"e�>��9!p�9�X�
�Uq��p8�!�nP,��텿&b���G�&�/7�Mt���D�*����=��j��ƫÒ|߫�4���'���ϫ"u�:iR$rcT~y5��[	QTZ���?��O����6.���X�(T���z���Z��u)ˏBc~RpBF$�RNUf�g�[�u��̸���������� �L�;�dD�Lg7�G
ǥ,�Y�������V��m᪞�{�R��W���GO����uo��g/k��.�ML2�[VZ2�o��#[�CT�[!!y�"����jF��dbt�s|n@@��Q7yGK3F����I?ѝ\�c)F3��S��g��[��P'T���g������H%c�{k����U�'$3]йw_M),�]8{��Ǟ�%�c}�{�^�)pJP"�Z�c����ɗB�ٛb��%	ڿ�wK���gT�A�vٻ��%��6DSǌ�
�w����MI;����M��I�q�u�$�톚	hK���|���N�	P��*λ�4�٧b�p��c� ���2�Z�!($lK�����?e��ݯ'�z�9%e�2���+��,RPN��us$��LS#�Ҡ[��,c(Z���~�dv���O�:DU���y�yV����
:I�	�%h���b�`{����w�����)�~έ��"e��C�Q���I)ܰ��b�ŝk��\�
��MXT^Z��-�t�2�i��EIl/A�4 ��T
�a	4;������6*C���ѱ)��&�¼�cT���j�Z*��Ҧ�
F'��\(+���F���*��t����A^�1���������Z�EW[P���>�(��|m��#9ߛ�2=��3�3(S���<��5H�L�f&~AJ�;A�����k�Z���"�|/��g��Nn��v�03f̶@`��7+�"�+���S�ﴛ���I������Cq���*v�喃z}��Lu���k��@��O[�1m��tpp����g�"o&_�{���.����M���n�Q��6�\.Lp;U�YZ��Ѓ���Nl����e�s:۰�~��aS����^����X6~�j��Q���Xۂ�I:W�i��2(5Lg�����?J�Q�)�g%��/Q}�M�5S�&fH\kG=7bu��F���k>u��>�:��y��o긺kld�����֪i��Iבּ��A�T���?��f���b*��#������P,�����	O/+�t���Aؠ�g��8��~pT.h&&��#`@F6�f��K��J;,��"��ɍiK�eX�U��)��$���&��W6��v�\B��Ey��/	Q���s�I3����m��Q^7�SuB@���v���됒�p`�Mh�cI�R�s��O��a$��蓣,�2~�o���=�9[��8u�7���ޫ��ʦ�sᾆ�4m���}��ߦ�4��yz
ײ;��vSǶ��b/D�}C�!�`Y�ey<�0^Z�A�hu�w�M(�����{2�����RcxA�@�Qк�u�Eo��Sy�s/olM�WW��bhj�_Y�?Y
ڻa}��pB��*�/���q�;nΙ�s������}��L���z�ϵP�M����]���ȋ�"RF����*ZK�j���΁"L]t6@}�#�Ϣh�^y�m�=�/���♿�P��M�`�X�k�p8筡�(��OO2>�z���8��"�W]Fr���m�6�7|ܗ��`9+Ohp�4U�0�~�M(��wC2�
F�x����m�e����l)*����E�>�E������W~��0J6�0�BM�<B������r>E2U���&U����O�3�?e��_Wl=f:·���#x�y-6Xa.<�屘�:/���9"9U�����DĲm�;�����\c�\h�YH%��'�uFr�t�:�����Z��۶�E�H$ x�ݨf濙�6�����p
�B �B��甕�(o*�����fG���0�Y ��b����'0���*l\�uxFP���J���M�xN�������U)H��8��bd� �?�����@Es*���XSb���5�O�&WSJ������R��D@��:�̀��2o���}���&c�|c�~3��&���釙#+oF��Z�m57�D�Nm2�N-:�!C��1i�6_�OE�s��g��"�9ɹ6F��j ������u��rx�.T$hc��l��r���"gK�HS�h˫T~l��n.�����F#�i�n��9��L'ڞn>�}�����l�ӫ-�6�*��Z�9�6�kY��j��O����d�q���1��+rĢ,U�l��s��,�H?tCX�F��Z�BX|Ov�Z�q��|��O���(lZ��n*2���y ��π����ymh �$l�[�lL��6�Y/�����Ѯ[DD���o�o�gY�D(i�&0�u6ܵaӊ�ǰ�8W�[כ�'^s�v�T�i��q�����ˀ6������O�D��D�����7�~c�t�"<��,>�P�T���<��p�#T�T0�������/U���I2'c�{� <�`���ˠ�ԷK����g	6Mg�CT_Fsj~�(G��C|1m ����6�e�^�����ؤ�'�"�*�ɗ�m�k�[�鑲F������n�]�~ڵ��Z�����S�����*q�BHYYh���2�����4�