��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)�K�7�jQѣC�5d<T�;Y��_'��W�!�ݾP��J�����|-�6��Jss�#�ic�	e�.�'�fh�q�1�w�	�O��ӑçcD��'�T�0$�G���.�y��8�ꁙ�KU�Hѽ]��͛;���\�נR�n1�H>�z!�LW�WY5q4��[P� �q�8a݇�a3��ǿ87�a��� �b��|�-�
�v�,0{�LIy�&~�NAa^GN��/d�H�˼B�8��'��&��t�L�J��\R$�D���0Q�֥�g���~v2_�Q"=�'������C�CD�M%��*/B�e���.{f���B��"�2�H�i;�����`��ُ��g[f���ji2og4��<D6a��x�Fr4����CC��֜3�魧%�㣻罴�s����"4�ߖ'@α��B��X�͎�BLM<Zg-�:W���[db;P�:��M�t����X8� �zb�c9O��`0w�[��G9�#b1G)��`C���)BXV�p��@�A��j��z��f�J �W�����NEE����j�6�Iޡ���h�}ʜ��_��D��^!މ=��n�&;��Z�I���W?��r1�זVP�w��V�u���莊;E!V���K���h��L��_���A\N$F�@�֯Ģ4�>�������}Vip��lc�zQC��~�HD���l�W�CP6­��^�����q�R��^��ч��F��O�ru��xF�Mho�W*�Z����'�������1	<T%�n嵬�#%�y�÷�8��BϿ���W���!�g !9{ҟh�8���QB�(�&�If)��J~l�n�E�����رVu0���"W=���j(�&���I������h���A;)�x��Z*���&��g��(�F �ӵ�ڿ-�?` ��|�ڗG�3a������O��8�\I��LVqR����P7?́ɧ'���2==E�e�=Qj�2E��b�����U�nuB�\/g'@c�箍��DMm���"�w���C�<��۪ �sRl�C��'5�����4i�ѝ�����oܐ�^�տY��. ���Yd�����~�f���L̨�pu"qw�W�i���C�w�b)M��E�K�TжiiN_v��ůw�U�������_cc�w=��a+k.�x� �܀w�[\��)�v=�?[�x -w��t_�����b J�zU��BO[�����(�?9U�����^aE�r�0@��aόF��7m��h.���)�DDJ�;��#���L��6C�T�Sج��Y!eL���w�ш�����c�^�q��f�A(�n�ҕm�I���8��C��w�h�j%�t��x_�'�//8�h�"��^Ojs���J�-�Xh���@+R�t�����ٍglYs���-\���.�7���o�!�4����t���<+��]�|�p�H����U��'ޗB�z���&W�R����n��^Z�T�F,<ն�s�@�tM��j�%�T��'r��-Bc	#����q��8��:G�L�u�b<��,R%~����n��m	�ܪ�_�>����\W*t��$DղV4K��#
�v�O����r�BT'�C*=x.�7+P6$�1\ց�����wz3�_H:����X�Ư�Z?�e^B��T8�Ž%8G6$�F�����ܟ߁H�-��*c�=�"?�AR"~{I~� |�]��\������h5q}KeC�w�9&J�ċ?��lFo$$6��<�$TT��.�nS���Upe�~��Y h.A>���,`5=��o�z���9���^�[V�_!vAE���e���0z�>^[do�JI���=�"D�4�E�mݪ�_nD�rݗ�v�U_���t;�a?�C����"���)f��.ܔ������8�Y�0�O$��_�	 D���'4/|�k����a�YuQ�|�jU��$�K4;R����V�@�BJ���q��\�K�[&%���Oǃ�U�G9g��ԙvƢ���3�@M��D��Mh�ل5���*1E��s�U6k��a�Ⲹ�Y�"��qf�f}Y�!O�U��AY�g异_��!:$��u���q	`�ig�/�3�iY�W��ȴ���(�v��,F�7��8c�� X����:��T�H(�P(����(�w�8/́$�#�G�B|BBR�l���y��"��|	S��E��\I���|$��A[�~ʓ�$uQHp>�����fG�6��k���zf.0��W��O�VX�ݖ���:Y[�:�Ǘ�d�����y��M��;�Xn/�< s�\l���q�kP�X����rPD��E��J��q�v��4
���ǅ���^�B��rK���iЋvj� Z�`{��	t	S.�R6rc����
�.ܫeF�HXЗ3���s�����M��*K��5�y�権�6��ݲz��NF��Lh�@7����9{~�.��񿍘1���8�oB5�j�\�� 3��:6eyvg0W�R0���2��d{�Ô���}�uH�.���b�r���*�Z����\a�X*8��J���]��/�7�2�Т�j�W�K��vQ��e�d+��o���솆- AU5㥇�:��ܙM�K oC���ɘZ���������#\$m駖0��!�.�|8c( 	z�;}V���a�;�Q&h��w0���Ǆ�=�ٺ�?��J߰g��>0E]�m4e�8.����ei�\`�2��>`�V�U����O�)o�AM�5
T� g��5���h	W{(�/�`�M��~��ơ$:�,~��TوV�4�H!� ��DU�n����w�sn��C,�`�z�y{��c�%���s�+@ڞ<f`�/���U���ͪt�p��]/�o��.�ȿ�Ȳ�A�"X��cv�a�@�2PN���:gԽ��N �f��@�?)1��W�&��w�jfԤty5���@���%,<!� 8�K͍��K�|������].�]~.s���������o��f�ƪ���11/V���{�x�Q�5�R�����@E������cM/Ӗ�p���q2Z�@�
7�(��+�6g��/���i�[���,�C׾]nBY��w	6��B�]��4H�����������r/f`��4����D.j��9<����N���&��tD���/c��FS��LwON�Go��	&�;��z݂��2��u
B��+s΂<Ѹ���.
n��E�0��D��Zh����Hh�9E���mS�6}݂l�"��w�+l�=	���n��Tx�}�-�?��5�gR�z�L=S�y�UݐBS#��r�b�@눈�RrJd�Ղ�Ɋ�5� ����8{�QW�n\l�h����=Re/H��x\��G��I�6��ECRo�y@C����lb| ����!x�b�ֱYnW�h)�(��&�0�X�i@ X�&N� �)Knj��F�jz�Jj�Ōb<�Т�ہ	���cq��"�Ui�K�&5k�{Y℅P� ��[ۚ/�|E�Qz�\��4��)7\�݊&��<j9?+�<n0�h��0~p�	�����[zɎ�˛�$�x����ү�����ӛ��},�� i>iF6*�^�GWw�P].P�b��ߩ�!@��k����I�C2��gN:B͐k"��T��Sy �����6�arY�q�@uS��֪g�a%n��\E��Tח�
�5^�dDG�<��6��}1�<���d�1�3h�u����SXT�N���2��M�tur�?(�Z�r� ��#��[s��#W/1�?2��.ֲ�\ ���Oq�"���(�z��T�8�L��&
�y���:��xwE=� e�9{C;rU��릃�I��'��̈́L^	J���y��ϫ#�@�%_լl1%B*d�bI]�O�j����r �D��)��1�.�H����4��<�H	������"�Ŧ��S���Q�k��R@�U�~�T��,������HĖ%:��-�ôb�>د6��%�X���1���AAEI�u��I��FFȐY���/6ڪ�M�Wz'���p��ޟ��]-M�o�"ȨV	�t���>+���P!��!	�>�wb��T�9�'�D�D�,�R�`��A��<KV���W��1Il�+'��3�؄�)��T��iJ�����!"V?Sh�
�V�Ń�7$�~��l�	��~�t��%�2�t��b�op�8��8�Џ��5�ш�� ,���	w�<\�uO���b� Hԣ����)�Tݺ��'H����N�A�0������Fh��\��g�?j��<�U��疝�o�3o�eAs�T��k�[K�%�h��䰺0��u�d�����av�bP*��R�3���gH8���?� ����l�3������Ru������潈
�R4gI@6���`K\�r^�懵��@J�#6
�_A9�[�5ȇB�+8�� qO-n@����6r�Zc�[K%�����j�.���qU7��!T�0 :. Y�f��QV�gLq�!�j{u�-����[�zby�f�@�f�6--�ɗ@�����n��`�~�q���������)x2����)+p��Rj�4�=
�Tj͘\SO��d�V�0���6ތ/Z �{��[��P`�%p!ڻ����d}���_�X��Υ��޶3r)ڡMR��?��w���;��:z����4	�ی��\���YW����>7��<���e���?�G�io& 	�uVz׬1|F	�sU�28�,~ˉ}���rL)U3`�x�|�T���.�#eb
������vA��G�����V���P�;��G;��ײ+P���y�|�ʼkR9�?��k�����t�|�-�4.Ȓrp_�{h�]2�b��ea���eL6�ܯ����:D���R5�=\���w PP�>�[x*��Ů��Nt;�D&����!@������D;��zy%�1��V̘^��\�NT�bi��g���*�G��l7��f�q�����ab���AȟRK���b��$�)��S���+/NV�n�XV��;>�wN.!�;�����2�[��B�P�'�_�*�@�Li�8�J����|h6����
��:�?_+L�C�X��$���3y��5d�NF���e�U*俯;>r��i)�&]�T{��_��#
[) �(��jfGy��� J��o�M��� �m+���s>]F��CR}��j1���8����Nq҈Y�����]�@&�<{��DO�9�����f�\Õ:kǧ�%�$�2��g����'�
��r7�w��l@93�-}	��T�ޫ���\��|�x���i��}���4\�?�Z1�Wl9 �.շ-X��L�Q���L����N��,����bq�^*A�U7q}��o|K��#������ �*1��F1+|�Q<WJ1n��j�5L�����jJr�y)����P����g��:1C4�A;���}-*馛{�t�Z�5E���������eb��H)��r��nV��9Xx"aࠫ�Ī�pӯ�o�Q�|!+O����Ce�L����x�w,�k�-�r�C�Q*�Jv�K��j�&;5G��U����h�#�jD��<�����XB�hd7�]:Ȟ�0o�P�P~DJjau���i4��a�+��r�Boehu+u���R$�%A���0\�ߒ���K
S�����3:�Q'��\�L�3�MY���8-��a�v�;?��~P�s��/���aCi���nN�R�;������]F��NW�]�3c%O1*�B �N�͋Q�h]��������o��t|�{!�
�.���Զj�+�W(�y�\;	�<9tɖLG*Щ�x#�X��m�w�&�������eG摴������ҟw��^{��
5.aU{f4=���~���������.~�����Li~j��?�S~W�j��~�]5�����߮���(K��û�A���	��0U�j�e���^����i"��V���H��q#!�X����՚�	@�!. Hl�U^c�m� l$���H��>�i�nʕC÷�ESɡ�pe6�"]�-���z���f��K�
��[�v�Z#X�� _хC����5�0���{Ps�����\� >���[�Iy0 ��y�qn�+ד�/_��eO�G�x���yv�F!�y�c�ҫ_�dgЪ�3s���Dk�=�\>��@R��V���Rq0����K����I�Kx��0����}i 
���3���B��<
C�6gvU��c�t`E��5�)�=%e�$Jv�}n�ͬ�s"�z�D����Ɨ9�
��>lfJ�wVzĝÉ��Tm��SO��J��r=i�k�H�A�C;���_Q�J�;��wh��ݣ`@��ƍ�	��
7T5��1v��0g��a	��I̤�d�y�I��F���G�)�f���a!�*��좣��l `~T3n�Ա�-e�~̚2M�#Q/�c�G�k���ϖU�}z��l�.���vF+���Um+��YV-q+���ʙ��#bUX�R�/��z.�~��^�ܲ�'/��{�#!	A^f�Sׄ	��w��ݟ�"��Y���P��ޝ3�q����=F�~l��(_o�_���'®�)���{�9�)���o$_*k�	L���* s��gc1,_� ���$7b�)�}A�H��7�z�����?QzQ4D��G,U;@��}-C����W�&�B`�J`�� �H�]9�r��(H�vƷM$�ܟ'wW9�M�iyXL��҄�|��%���SYC��I�AtOқ���÷��-�<� `�������:}�(h�6]O�ة�N�ϮW儱�3�57C�mơ��i�?�������f���~Iq���ַ�o��4m8����o��C���KW��HdE��&7Y����B@��E�7���ϱ¶�z��f!��>�Lњ����r�=پP	�mIߨ��DZ0.l�A�^3ԏp����f�NY}������\QWj[�KАl�B�r���rW3T�1�}p���8��L'�V��'.)Ȋ��\4F���,aӱ����23?:?��FP�-kG�7�$����._,rJ�0Ц�@�
1J�y�n��f�]�H���P� �~���#֖��k��A��v�Ʒ+��b�$��1�o�M�)N1Rq�!�h��~�+<U�s�Á�� 1o'z"뉥�p+N�t�;�p��Ԑ��o@�E�HK�7:�r2��Y���c�� v��y�z�A�T���¥8�T�7�r���@PG�}E�ﲘ�ج��6���ѩjN�k/;�j�v�c��L����GL�F�[��w��^w��p~Q���s斔[������ ��`�˂�=���M�\PUA�݌��G]�4oM����^�P6��fLqB"��w76OKi<'���g�V:�U�5dס�^Hl�CY0�H��aB�mK�-�d4�Շ�BTN���8G�8����[˽_�LZ�����A�Y
�2t����ÅM�=���b��ԭ��~��'9D�d��h!_��^5�VW Ɲ%)w�5����Fy^Jf���5�" ��(ä�\��"��>��iFxT:>��!�d�(`��|3��o �"�A\T��m�P�r��Q�1=m�B1�bs�4�F�x"a�����F�˦��N�0�s���4�4��!~���֤L'����	^�@�ґ�3��̊�n�0LkPT{c�H�V��Fy�����j
������Æg$O����|s��P��=���v�txk�+n�ewLku����������)7`�#���K�z6�JTܒ���,��N�7*\5�c�����@j����'��c-9<[p��q҉5��M5A=m*�kt�T�%z�z섂O
+ ≏a�od{���(����|�{?,�M�ѵN���ӯ5��� a$��HS�@o�����P���o=m����Z�W8�4�|��c�uB��o�Fo�[�>�i���A����}�0v��[ ^gx�8�iV>��ģ󾶯�T=k�ڼ|���W}Ɵl�'������&�G���L�r۰��8Ҙ�>
M�tV"o��z!"V�>�Zm��7)}�
�&R�Q�C�\��i=���?�"�"ïo�B�	lB_��k��N;��Jb�;�L~�X3a�k�C��{QHJԝ�;�9��zfSx�t�ʵ2�wPq�/30Ջ1*\D�L�?q�:��T���^3+xCA�6`������&�B��Ҭ��+�|K�/)�h�@؇eq/0�;WV�q���lT�׸�X�t�ݏ����OVG��\��"x���Z��۾;�.�ǣuO��0g�Q�}�o*������t�����}E����0;�A�C��M��\}��a� ���b���޻Lw����ˮ�ǻ�q;Ga���l�X�8b�Z6�⑯t�m��"O����[��
h�c�c�?^`�H��i�<y��.g���eN��XL"Fؖ5�ҋ���iyG1�Z0��{��iqmu`�D�{��kT��E��U�_W:Pa����(�V%�'�{O��q��E�u%<�l)�
Elx� ��4�xq�,���� �3D�������OwX͋~іr��:t
���h�]��$���<�? ��ï}���&�J��Zh��!��ZA8\�5X �eO�^�C>Ӕqn����/�S�2q��)�J؁*f�x��D��Z���h;�u�(���@����yl������� +�e07��l�%n�����9K��鯽5��L��i��eH�:{|Ġ'����D@ �x:3עe�,�D��h�z�k/�E�Q��+���iy�	�M�x���V1��Ū�'1�w���Ve&4�߽�s3����i�OF{_!��_�۰;%�]�sλ���K�}�1Q�`�ۨ�p�`o�����}�L83[�`��v�A�սJ�_�TJ0�*��
U	��1y�v*)tC���tXXP�*�)���}FY�,�+O����@�|��PП��� G�wv�@u���i;���(�����3]����Y���"]��膢I�b")-�y�@�6���8�S�	\b�����	�K�߸i��*�gɐ�ٍ91� �F�j�s?��9��aΏL����~=J�ר�F:G���q���7�uQ%
!�	7��P�w�5{$�.��b�N�*o�?��!Z��N��c��Q�o97+�>
��C1�;����b�qa�(8���9�!ӱ�m%�o����IX�Y(3�J��;�ʁ'PK5�xL����f\c#O)f?�N^�r�.K�����R�/�w*���B¤R��L2������S`�i�v>�B�'�����
�ڜ)���#�~α�ctJE�n[�#ݷ�we��nP'�XZ�8�H]MP���̎�*�G�x�\~Z'��
�G5�����i��s[��k�9Pī]X��<�i��y=�
k#��i��6�vܜ
��t��C��a�s�~����P��;��o�Qݕ�D8���{��篟X�;��g��gt�f:��,�g^!��H��3���I��>���:n�i٣S=៕�Pq�+V͵���Ǟ���h�EF懁O�7���brt�����w��ێ5N��[(I�4��^��r^��:'�	*&�G6�9u:�ye>_@Ƿ&@v{L�"���<�z&���l�
	�H�i��.V�����}Ş�V��2��kD�,�}i>oU�}�D�t�,<$G"b�\j��ջ�؟ ��!5 )X�hڜʎ���}|ZRR�G�XJ̊�&9��OrK��'̝�޽0�Ԯ��%"H� ��^_|L��e�9"�գ�Re��0g
�x� ��u����U�H��������)�9u�`��*HL)��g���oL�Ǧ�T������X�,�Ug������I͛\I�VnX�w�38�����a�>��i������T�&���Ƙ��kWQ��7�lJ�aR�n���Կ���B�ե� �����&��{b<ʹdRH+�/�L��P���Ɵ�Aa{���;�O3mr,�v��z߭��â4���7黻��)8of�2����s�Ip�[9-n�|~	��G�`�5�_*�?4YQ OC��3��Ѯ��_N�!�-f����N��Ư1gb}N�)^�o�`R��*�w{e�[�.�M�n�r��T5U<S3�
����AZ�N�Jg��P`n�P�J���G�R�]�?8vL��G��#�fz�n��&��݅��:�B%nDgd�X�i,��R����n��3�n�a��j�Z����"pܺRVd�}`�(�����w��}����7�k����^�
��c!����0�Vq��k�ً�Z6 !w�K�ACKÜL�7_�<��<�&����ޭi=r����t�@������Jm�E����@�O�l]�ӑ���Q�l�ze�;N���N>8�k���5;ۡGl����5�mk��!�5�E�;���5���8{\���u��0�?4�����IR�F>#�5v]H�[d���:e� ��r����0�
�n;0���%�ry�ƨEm�*�ϟ�ώ1���@�V���3��X�uʍ*`���L.��.���!zV�W�{���I��!�F�j�8i���:�W�5\�h.8j���O����sw/��"ga+�X��l$5�~P��9)��n|�#���pO1�k�é��vs>�7:��nqNL4�H�e~Zx��C黠������/�{��$�(��\� ����/�]�����uL����h��k��t[Yu���<?=��L�FiS3�)��{���e�S�2�BEjuz<�B{�A��듇�n��3[d���|d���_��`f/�+��z��>���%��8Rvan��c�����e�[CV1/�k���U�x��k��������
Y�#fZ�0��@��!�J�C��S8H��45�����lx\�������"2ƕ�S����t�z��l�TB�%v��2�4���{F3⩬<@�R�/,�gu��b����-�?l@�L��r���ZQw�]I�ɡ2�k�S����/N�a�Z���ʒ9�e2�	
�� 1���*���s��c����8�
¶aʩb݊@��?�0��s�Gi�d�BB�YҰ�X��
�ӆ4��y?�m�O���y�����݁D�+������ݚA���p�u7*�~7�BWi��<'#�'�*P
��ir��clR��������P	މ"�mt����VX��S��|�\��bɱ]��� jT��ݷ-�T �B/�=5J��O��_��.�]/�\z)i���-��������=�<��	z��R�Ч��,4{�ֱݪ|	�#� �H�|+�`3�[)I�85�	�v-]#���37O@R���1�(G�M�O�j߀ 9u��Y�l�S
�~}<���	Ѣ!�[������9�
�3�A}v��s����O���:�b����n�q#��U�'�Q���$B&s�`;����
�"e���E�Ό<��'Fb#Ñ1�T7Qq�'.��M)��Z���+���+ۥ�w��^���4A�!�0l�«���?b�u�����ec�u�TL�$�=��G�A)��0atK���
�ޅ�~��X>�0�Yj��z{*���G8���qB�ׇ��̑o*#FO���Ǩt��wm���y��6��<��Ur��(�+�@
T�C�2�E�f���T$��+T>e]!�#o:�i�B}e
�����g���H�,2b��R�NsF�x/9�<84��V���H�L��;r���/w-7���k��h�|@<��^��a�ށ�	�;���M�gb	jnsw@l��"�v�0���&h���m�I�3��yEg*e�{j�=元ȱ�$j,h�e��O�Nu�&'ywEt�5�a�`O���s/3<7<y�Uk�u�X��xmr�Nʚ&�����+Q1RjrPeܙo��y��	��C������d��^��q{@}�B~\�m�ú����q����5,.�Ңp�d��PH�Ab��~W�M����U��:���<p����
zD�iU�_]����g�$�EJ	�Urϧ���iY�!�-�l�&N���R�S��n����������A��LVcM9qV����:C�l�+�������.�m�Q��|vF#e!�L����١d13�M�#'�����T]&�K�Vy1�S���Q%�;��q�!�uK��/�$nZ��d��d�ne�i�[�t��=��4l�\��]��k/��qpkY�1��ͨXz�e�rv�Q��Sj�g�˅�Xr"@�3]迧�.�~8�����َ$g��$�<Js��U�]g��;j�
Ŕ �YZ��~z|� �b��v8Y}��<����:��?9�d�Hn��5�|C�}6_�jU���{ w��S��/��"?F��dDB���?��l&�JY0:�V�7�:L0&���o"X�ix��a֘>�3`��$���x���9�� �ե�G�i��\�3+�~�>SB-���?,]�H�%�NK(]l���3�"B��|s����~Bz�rބ�'<W��W,0Gu�W4P}S)�?���|v�w:X�C􁮪,>t޸�}���L���>��119���&��	7��R������eY72���a����yk���ݒ��~��S�4r=*�\(�y�5��QO3�tiy���t*��Ӽ��+6АJ8t��m���RTg�ʳ����Y/{�1�)O�$���7��
-�P�H�wʠ��2>���;,��h>���V����h��X�s�I�H�<Ŭ6.�2��W!]9H�]��v�.g%�q��l+����쯭0��4�˂<���E����N���[����y�T��q�{΀�F�n�z* u^�ڝ��1��Ook4�蝖'O
Xe��G��\i
(��R&&�E����:��M5�٪Rly$F�#8?�2��H/����vd��僸�v��;k�.H]���(J@#�ɘ����˘>�`F W �������N�M�{�%v�A�J)��4e��w��ZCWy����IW�{%�&3#�N���S━�+�a[l��+�x5�0�Հ�h���㾲����`�rX�ŏ	zԎZ#�\<t�xZ�W>lXX�����0��W3�O�F�BD���n,]E|���Ѐ b��,�c��FTug�`3�|��<T���Wջo�b�_h���i�=CK�pBk�s�b\�� ���p<My��<��sl���,�$�B�!�a�b'������M
Gː��`փ(��ed/�p��9;��U��;Xc�[�<&-A3Tk��fŻ(�7(S���#�
ԟW����!�)��x��a7P�?�w{��'.U��ų��J�$a!��Y���d���t#�S�^W�D�Vg�G�Eg��z��<����oafϖ3I�ti���$�Ֆ���W,�	+$��'�'y�HQ��������D�Gvjs�qu �K�����xN:Ҭ�g��3��uǿ��D�Ұpދ�
uҒ��x�H����I�1s���Y�f3\����jű�"\@t�D_>�2u�f�#�oI�n���)����C���9�|#0��/��I#��?P�hn���K++9�1���X��A<��Z����׹�H����e�ʗ���P1�pk64�%l�e���i���p?�~0����>�iF*���g�'�-���h�N��t�̃9�2�
��G/wS�/�3�3�\;��bF�8���iJ $q�ʏg���֠9.�K&�T�L.�Y����÷R ��7)�3}�l�������)䛓D#�S���Pʆ5�~�p	;$5���/	\�	��^����?է�$@�i�nU���8�H�M8��(��H�,+}�?KI���C5��N/s+Q,��2�u���k�e�$�U7����E��]��V�N"ID��$�E^x�)�t��
"�Q�j�h��a�VI�]��bq�o;��T��
0癨�Ƶ>�9�T��F��.r�e���㞥>�e�-ē�]�X�Pw���сU�e"���s0c���Y��co]�CW�ğF��}�ʣK5��+P�=f��:7�<�o��YD.�p{(�#�
u��������;�-M^�M=�ŔM�)	��)��(`XEs��z~���o���wn��){�Ʉ�f�t-ᮾY6�0c2������X��Zb¥|���Vf.���462�g�8��Η�Ńy"4~�ۑݲx�Bb�A3	�Drz�\�a��Z)�����%��2͊��v�15"��~�v��nұ��ׄ�(: `?�#��!�m}��_Fy�1�@�`�ր�L$5����3��U���c�B�jK��UOإW!�t�#��\��M��J�[��V��3{](���+ɽ��(����5e#f�TT��ȫ�[�7����Q��f�e�g���2�j�l����p�&���e��nbr�2�*߁<�G��JŦD��l��&\axe�eR�T��GK�%h��S�j�˓��HH��Q 1AI�ux�[W�;�c�U��?�p�ߩ�)����R�2(��,��9���=d��0�16����X�^�
e�{��A���Z��0�0��0�n%���H�-�����rd	ˍD�m��3��7d��d[D���6bn�0�<{"" �}s�9��1*5m��a&������֛eZY�K��cg5.S_`*��J�y�q1�'#t����̘(�KP�lN��7|l/��
b%p,��u9�~�iN5��L������Z�o�a*�S�hP%��\���l{���;xu�6��\���88�����$L10�vo�n�깱�px�4�,�m񃊫P��!(u�ire2���]����aC,zܬ�	p�V{\J3T�A�����HT,�z�L��),N}��7��2r)�H��whf��}RI�[��'������.��˦5C�}d<	w�x<��\���w�E
��^�3��#�D/�uć��c��;�@,�5���	ʹ���N	��O��m�M��_�pb~	�s��}�c�|� �&!��L����3���睍@^r)x��PP�s�P9����B� z�����,�L��ë�ñ����O.�ooGKlgҸ����çE���luM�=��/4{�N����5 8�7Q�[Щ7�A�Vo��wc�t�\yKq�
��ꌸ���Vd��P�B8�N���)�;<��bk�Τ�vsf�әWٜ_U�k�E�K%�s�t��u ZD5��D��l�l���F�.��iM4G�[q͹���.'x�w3��
�bh�463K)�����l�{���o�<S�DV�jo�4�w����;�-Ё%h��^�P���~����f9Eɸ�]���a�.W��&u/i�'Jj�y�N&ZtcG�-ߔ�4�[����T�!7��o��w�Ӏ����񅐴�	�/h��DșϠ{y@4�WY�A�*K3����`�kFxk��w�6��� �����22��f�9�A�%<��'��v��0� �����LD0$���f@�	��M�q��4�9D���,�,�#ȍ�(�VKŪ.����a��r�&"���"Ѿ}��M1����X��aCe:�Y�����A�?�ɠ�lg��p��t�.����d�XJ��̬�����Q��q*�'�#IC"��,���nr�Q�+U������I��`��9��7�U�}��x�	�Z x��K}�A�,z�&�e,㭜���\�j!O�v���Cow:�����Qw��o������'þD?���e\Bo� ���>x�F��d=��@/����@��v(��*<5�a��9VJ���I�nx7�#����_[�����ms\���?ړ��ݏ��t���*~O� ����~�ir	n6Ey��	谿R�	���9��x>�-B�g3�����H� ���+Y�IWs�k0�9���#��wr�9뾢w���5����J���C���8�)�#IJ����P��c����y�ND�9�T��N_�W[g���١H8�����Ay6�`P�ۙ�����\*q�݈�Nʂ�2	gu1-ݙ�gz�r�g��T@P� <YF��%pRD�W�_���F6�nb���L��лE���IYE����WƂBfI^���!Ҷy¯�j�):K]��ٺ��v RFȦ���$���]�F�`�D^,�����1��8|	;�z�Pc������o��1��H7q��U�� r����"dH2y2�z�ُ��
�}�P��,NP��V��wo����Z�&<�za~w��~cy��-ʝ7_����'d�D0�!8ze;�6)[����0�����,�
Q~�̅����[���<(��I��`��Q������EC�D$ʉS��f)�N��zEo6Ѳ�7�� �4"A"�^�˯��X�9���|t���S�M�,�Y%��@��_����-6��Y4@(���l�����~�2c�v��n��h��Qvi�_�y��kD¦V��Z�w;:�b �m1&�&{wm��?<>��k�f��%�s>�.�Z��+���\�� �>������ij�еi���6Fga�ƶKF�ժj5�>�kޭ���H��IdS�E+��Ԉ�7u=w丶����*��3ʗ���}���,��"^`0K����wIu���U�YM��+ڿ�����b��4@�sꀪLH�tm��7/�J�G�VO���*$a~��b؈�7��Ϥ��l�rQG� #y��n\����f찹����io���{w�	�v�	���)�c� .���@�f� q&�A}b��?w(�3�U�K�`��h␪�7DΖ�#�+��� z_��z��7���1�	��G��A��s��U*��р�a\Ɯ��4y9�s��������Ծ�-%t�Ӫ�WB�{RW�#PrQT�9�7���@39�'��ZT���c��`i�p&����#w�Ʌx�eF�;\yDU��Xe?h;� PK�nV�ꖥ���]g����
Q8-�mz縡+$w�X�>`U�0!]\�88�x<؍Uw���_>�ŧ<�ɣy����t�q����Ptp���n{k�+�'�����<M��r/)�#�?��<�~�^���%��<��l
m��a?�IVz4�FxVy��֝�9���P�_��v��o�R��)ݍ%M�9�i��h��oΉ�i�H҅�j�)��^�1!lm�e�1֝vӎ@�mN�Ђ�D��,�E���4�s��~�L�(�0��SH!���\5���Á���@D�n�o�;�L�����j���s����թ��K��3�c�����@�pC�ŧ��`&����k��r�c0+���
+��ͣ#�������M�B�rmD�S;��4ŖPc��G��󨐣V��'�{ރ�|H�􅧊�E'��}��:�<%Rp/��Ŕys`܋��Q~��u=��Ԩ���zx�O~�`�6�`C��ܐ��WW]OddE���,dj˂�bn�y�_�{� ���A�3Ю�d\��-a�_���!�Z������ie�ԗ��`�7pn#z�(�a���ǋ܅�W��\�'tڞG�Z�Sj+P��N��̋�£����O�j�m�
Qo�3��Je�x���Y���+zƶ?�������)���l�`����Y�:G���>x%%ath	w)�J��1%+���M[1+����]�
+H�dzWǚe�#7�ثg��D�<c-�9_$�K3�����MRv��[c�R��q�W[�"���`稄(�K|]ᤩxC+���ve�X�����w���ܧ�o�<_H�A�oŬ�/���t�9@� �؄�fp�P1��C��Z����2<�{�bcD*��iUO�4�ƣ��XЉ&F�ϋ�(6ϊg�|��hӔ���^�Y����	1R~��+�R)p#��P������3ǜ�0�%�x�?s�d�D�d�^.�JĬnb���M�'6<�_�wL�7�G��	/��7��ğJ�p���� �J�P�C��z 7���G(��ҥ"@$�-��K`D����.��1Q"�v�v:��
���^��U9�<�h
a����'������Lǋ��ADBmp���"	#��f`�U�Us�F-��y��F�U�i�a�'b"_�����0Ei�$����'mzOLNQc>8>����H�^#	]ʱ;��F�Zym]�����t��6�O���1-(��;���F��|�e�||Y[``�o�S������c�@��ά��&y�)���_~8��l�;�һl����PSK��HQ|��1��O޳�����
-�����6���z��V%�vn�GјW��.T�7C폖���k�ې�r���8��W�0�c�)z��\�����z�I_�*��I`A��/��^Z� �v++|����'�^����׼�0xy��7���LָW�K_��}r�e�v�g�����'?J�?�z.�P�ח��/����
��a8GV07f�%��A�@���(�o�C�YT�Ve�D��SF�~�E�̥3Cc5�^��<
zgQ'�)<��VB�/g3@ݧ�Y��_�Oa���}�d�teX#"׭P�n6����c��q@a`�6��NZ��Q�ĦBq�C�Gd#�宔:�i��)���NXi5m�����B8�����a��LӢ������
з:ߎ
g^��jOt�Ī��!�)�"�'�I�Bumuc'$�į���R|�j���J��'}�I3`tC��E�,��$�����#{�}���<kz��=�E�j�9Y��,q
��A�U�^-����d���6' #農����2��BF����
�*c�x��Ǉ�!E�xc����U�=⡅��Y�HG4B"U�'��U���3@�mfV�u��Fa�QMa�Fxh��6��c�m��@k싶���;TGى�\�)R�=��Q�� p賯�]t�K�У\d�䬳�\�j��������^�0� @���\AٗR	���mP��!U;���`���|��e	:/��[�{|	�#��R��a��&�1a�9
T� �Nܑ�B�p��]G�i։O��O�	?ak�����0j�~ȗ)t�m��P���}� u$��>�>1����/�=�B��9�C3�����*+���^o�s�'c��"D"%�?�>�)S�Zx5/y��r�ɶS��b�ٱ;��5�t,����W/��f/���e�}��;��Y�;{?<�j���/Ԍ���f�TBH\UZ���i���U��Y�pf5���H���g�<�b�S���/����E�j`r�zj�1_We��A������NT'$����[��.�;�H�����.�0�v֝]Uud�U����+�ݪ�?r{V��kf#���N!L��̽��u�-ԛ�^����׾��`�|]]`	T����YxD�,���c�&�Frh�_�҆/�4Ha OT�z�Ű��2.�o��?�������=��:����Y#$��8���U�����
d���(�GE����@.QrYv���((8\��w�(�6BG��g���ܐ龉�`�z�,����9�9=Qܛɸ</�/��g���H)huN��$�.FW��TM�n�.DMQt�YzM�Z��ɕ���?�>�wmL�����6o�ǛPv����)�������܋��^�� �}?�)�yΌ=pa ��c@J���n� ۵�gA�Tc��т*2D
!������徺Z�O�'��f��t�2g�@����� lf����#���Y����\�n#��Og9�0S1}���Fz[zV���>��ޅ����!�5}�\
\���O�m;���u��Y�6��e�w��KI� a
��6ٍ�j)׎+}�l�Dҿ��g��?���N����F�,���x&[ÝG8�����@YЬ=}Y$�@��Z�i@��Ŕi#�oR՜����̘��i�P��.��*�r���6q�A��������)��Q�@ԓm�|˨Ŀ����nF�ſ� &:��)8��S"��2#P&������e��Ae-�\-��;Gt�?Mm�����&pM�x�~�K���_����qۜ�u�9t�w`яXX�<�WX��p܀
ҐRx��ŇP��Q�aF2�W���KQʦח<q'5�+$7~w�2�.�k�krh��P߰7W)�키I��=�& ��ث�C�p�\�5��%Y�����hRI�S�C�ƥ�k��z�hG�1��XL�'R\�۵|����f��p�Ik����-bߐ�l^�T�D�x������MJ׾�V�4Y�>C�#_�i/��2x���c���}���E��CJ{��g�#�����C��p�b�3���-˸��gG�f����^�'�
KO���EϰKEқ��Or�����!kI�A}@�d������5��oU��oEy�D����lr<E��ɐ�����Kv85+O^��y?�ԩ��4���o�W��W�͖�ؗ|afb�ǘ>^�I"K�?���O= n
Mp���rO
����:%x����^���,�%�~�%O���͍Io#�7cI������h�E������N�%��ϻ��W�Unb:"DE��/�A*�谴%��ٱ��㋨�C�^ 59�<��",�С��"E2�����c�_���E;��~�W�`�Z<�@M�o��>J9<�+�)�x�y>_�����3�Ʋ605tpk6͛W�7��P\��:��C�?~p����J��@_�u�Ć@p'"TȈ��ߠ�~���"�*��OAz�37Nf^��r�l�* hdI��#	�x:��*�R2�gf2WaĖaֱ��]�G�*00zD)���{����|[��y�>�W��a��)w�z�7��%�Ћ������U�Ѳ��I�ↄ�Q�&>�yi���z#���f��;{����=�(	ejd/���Yo�o���S |Y��Y̏0-�}�N�F?f����p0q�+Kl\��߃�.���F�V�PP�%uR�\�#���"�um������B��ؔ8�Z�T)f���y���"ǟ�<G��z뻧��f� E�����Z��b�c�H����%�m�JolB@��5V���۱��H�S������qI�/I�{��\N��.���$/�tJV!�L��#}�;l��A�d*�ؕ#K^���%/�}s��E��=Ij����g�kr$de���H��Pw'>N�7)!�?�@^�I�綪��W�c�xa�n��J]�Kb��Yf�9C�Cp�ς2�7��� �[�
&@s����V��[��t�uL�%�&*q\��*�����|�ڕ�[�����R*t�a�v9%�]Z/'9�`�3���DF_|���i��W�Z���FZmLNR�U��[X��`��$k�4e$ХO��]��p�@~�vP�:�>����U����'���86�֌c�(Ƹ����y�a�>�O�t���J1����D�1�q�v�@�B�#I!��Ւ�����x�4��v���Lj�[����(��=DU���L�
����:�P��g�Q��Q���i��*����g��}���ĺ�2ro�'��&���d��ve�4���?]r
D@��N;�  b��iK?ȥ��af/���U��B��}�"�1_�d���0�/��-Q�S�Ku{����=�j~l�WxW�\�,��pV}F�5��_�Ϫ7E�� Tj'F��vs�ެx^ZOT>��r���q���Q��ͬpzn̯��ߣ;�r�m�
�f��39<"�}���[�G�bp�Ꮿ/݃�>�1�b��~�!"��+�=&ݹ��=�Mݸ�V����B3(�`�D!P��U8�H.hd	"\�!%m�^dC/Rٜw�an�1TTn'�9y�J,("�F�� ��׬W)��oȉ�3=̙Ź".AW�e��n�og5M�P
��>���U _�qs�hm��؞�=!܄}�6YD��g�>|�q�E�fFKd�W�V0�'vB�~?��q|�?8嘽���#)�u%pI�tDe{�/������o�oHO~�.I����s�8 K��'�|%�4φ���deo�_��,�'�kV�*���[�-�\%�N>�F�e���l v
/�>s�3��*T � �A<�X o�-�[Gl�p#W��YzLjhg�#wf:4x�1�b�@.}�`����+�x�1��:9޳�L�$W���M�M���a�@�c�Z�*Sl�&&D1ۀ-�;Y�UHx}�P��J'��X����k���Y+ <���)��=ǻ�����7����;����#������:����^�3GE\���dR8�,�:��	guع�a�m����姢�nP�g���zz�>�n���c�@� �m���*�&�=�?���
)�F⺉�~^_o[��5�W("_���P�����<��h���Y�F`%�p,	Z�}����4-ﯓ%�c����<km�0��8�E$��#�Z������w�(p��b�ޕC���1��p;!0[Ǡ��Z;$�8�Rj2I���<��+��+�����f{�i��}���<���;0�x���W&`ׇW�T�:+�Gm\E(Ť��O���ώ���U�+#�Py��<�k�@n�i�o���萾/PP�e�Vt�1��X��(�H� �0�X�y�nX��C�[Rc���6��p��Lۀ�Ñ�����	�_qjG39��-dx�c���o��c�>.����0J�#���m��C�\����%��Pؓwa�8m���Ku�|j�d�1�]��%���A��3�4���$����&V�
��g�W�D#��Ӏ�@��K���m�D��"�(�0��c����Bq7I���V���c8�lۈ�d�9ﺠ��fj;Za�2~��x�{����J�^�w���&aZΘ�BuQ��>{ ǧO��x��)�|�W�|i��O�9�Ϭ�Z�_pd���P%GS'���ŕPn���&�0��a��	a9h�Ӹ����K����F!yK&�Z�F��'N�+�~�� I9���yJ(�3g��;�f�-�� �.d"Ll90t��%7~�203�̦��>����G�3��L�������}�3s��r������J��XM	Ќ����G��	�V�5h/C��6'�W�~W�bX��@P6�u�d;���_X�rI1ˀ�*t������v�,�^E���qY`��hH��}Թ���
�