��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��I�v�aНҫr��@��oe�5=[#��r~J�z�v�HA/�\�xI�Ь�1�_W�t��~�~�ܙ��s�w���z�{0Y�9g/:�!�$����A�y/w]x;��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2���Z[@yh�̟3C����Q<���d��lS[�z�n���������F'��E�w.�Zv&���2�7�f�K�m�}��_tsgz���Q��r$H�+���<ޤ�I��;6�g;��y��P��I�A��:o=�5X�+��t��7�| C�@]�z)Bpa������d�d_��79�*[��E�؀�'���+1~ᮕEj5c������3���*/,q�{s� B��80NJ�W��������#w�BS�O����1�:�MS��ˮޢQ�r��/v^��y�9�Tp#Ƌd^�V���ڔ�ouq��P)���*p���+��B�p99��5� �j��i���0�a���"���Y<���p����<y�۟/OXa��i]�ZBL�
���qg2\NS$�$॰�ؙ%	�`*�D��;@]o��ו�/Гۍ����-�#0�`ii��B����D�
�����cv��w1���
v�]�K�6k�4���im�H� u|�붔Dm6��{��o���K/ yG�T����4�ŗГs��D;+���Ņ��D��O���d�Ô���qXe)�2������2p|�t����9)|����M����~���Y��ig!�h2�8Ǵ-�?��TnO��i�!Y�� "7�jl*�>�n,���Z8�D��]S��M|ʡ�4��9B+��U�N�J�q�[\��f��F��qx%e�K�����^�;�0�s�u��w^OrZ8w� I:�M[Ɉg���+�Ь�����*�y��
��l�;�AC�UnK�����
C1� �`(��Nom�4:w��jҥ&����{��;y����F����uხ�f�{��UC��xf�FgQ��(L�������'N�>N����1��[�d�c�d��XP�eE�.�ۗ��cV�uzKQ&�5��ԩ�~��yo�N�8�<U�򫖘��5��+��U�����j;���'}��\���} �'�V�4�R��y��0�~wHG��"�>�f/�)(�P���=�����B����-�����	�N�<�U�Qp�D8��^ǐ)׃�փ6���:��Z5 �4��^<�hre�ᦒ�j�j�s8��"m�%�ƆFF�.�$��	�t�R��yG��Qn�f����`Q�o�� �S�fR�H�D��=�@�b�#�H˾R1�he�@)U/Z�W#���.��l�y�:ʶ]��X��x��G�����}��f݅�@=������J���v��)h��D^��2(�s�I��3�῟���kCF@pp�e/� K��w<�zW��A�駋�U��a�ܿ3F�!�-��'\�w��[li�� �qֺ����8�S���r^��W|��2m xs��	��AiJ�l�W2��1ij7���Z��L��*�a�Vm��%��V�Y�eL���q&��7L������5� Υ>(V���q?���B�v�m)���Dr	�7m�K�~�"��uK���WͰ�?d�W��5��|΃xsC�sY�6����b濭�s�\�.3�����v�}�#�s���+����L*�T�n�lLрsi�MdB�˲^��x��{�{��B �S��P&>w��Ձ"<����~��n��9,y�@��=������<�4�{�C����9X"�I���Lk#��P�� ����+�?Edy|��d�Pq�_��
w�^ݞ��Mk� ����zu֔14^[1�-����^���1�#�C@�6��8�O�"�c��vPV�8\��;1�@�h5)��MM�������?<ުK\)Ь�&�������gBo������-��glf��3+�9�U	���0]�!|c�$8��._�� K� �6���0�Y�vv�1���1��X$��X����Ջ�v���EkA�xڏ��j8X<
�/W3�WDy��u��Ȩm��8YpU�k�F��a�(#��7����i~�\�3=�d0��V5'��mՁ���4mS|�Ȭ�"��7\�ӷc��ä5�������E�����X��Ҿ4�:�G�M,��b��!����íz�\�5������|?l�����~ƫ��W�Y�l7wן�f���*#��U/��5����b���H������<_*b.��b��4 (��d��诤h^�0<m˩��0�T�(�4����Vg�����yq��t̬J���|6��ɦr���7mx���CB�9ܚ�^J�Jľl��b���l(��BA=KDƔ�{#�����5P�dcP��w�v�Z��a�����A#�V�{��c8{�5�{�]Y�D���ag
�q���9�H���j"��* �or60���O�hȭ&g��;=�C��G| ����
B������]�0BZ�.pJ�4���,�/�d�>�4�R���'�x��6�𯽩=�����|��}�S�R�ig�
�{�c�r}<y�X�F�&�o���k�,U\�2�~Zލ�'X�"a�� I��w9.a�A�dwe�<�`��.�/qڗ6mni�bp6��+��P���K[�J�$v�ܢ[|[?$�51@��Acv�]s	Cu��.��#�s���p�4tS���ϟ��Iѵ_�m컸��a�I
��C���[L��̸\c��?v�o�z�c�x{�X�&�JZi�ż���':�@��h�s(?�~ë=�r��x�4�[�G	�E|`"��I~�Ů�R��'d�z�@��4�$I{�yڇV� 5��r��l����
����D��~���"w��FI�|gt�e�qO���a����d5�x8.X&'PV���c�������'��ج ���͒��\�)��Z�������̸�5�X�W��h����4��G�r��+�ґ/tTr��l�ec�:��[��'��Kj�^��ӝ*���[��*^ݷ"e�Y^AU^`����󪹍��@O���3U���쩕��3�ӠM��[���Kp�X�r��W	p��̏f�K t"�-6,+��c���.ǍI(����I&�j撓�R�!j�"�7�ߝa\�� d���8�5��!QY�JBi@�j�08��޴2\x�'Q?u����od�����>���A��8:�N�m" m�	Iv��8H��"���!�9�����+T��cl�hu�����CkD��H�_X����#M�5˖�����b�ِ�#��*��Q��)�,Q������]�7�Dv�b<�>qG�'hd�
����Х+�p������lAo�X���s-�(�3vuD4%"D���l�£enCc�m/�I8��Iwh�_���6'�%��H!I��#���s �n`�Ӻv��:�4"��>�
u$�F]�VT
�r�Г[�̊�ߟH� 
Z��6�n��ǭ�eV���&��5�	o1o)�rsc4@�WL��-&��jSP���EZ��9G�ř�����
�뇓G�lr(F�DGxM�Gʢ���1@%�?LqL��ȕg�MƎ-�Z��C,f6���P�(X.I�������dz�3u�ku1�vD���������y��f� ��>M��M�Kz��Uc�LX ��p?7�D��h���Ğ%5�EG�����$f>i!�rڢ^e�J��O�m�S��[
������$��������U��'����".��k�����)��E����p�h��hx��D��k}�,�LE�}
���,0R��@l��`k�K�%r��ܟ�D�P�����c"�F:�x�(:΋9Nh� ���ѓ���iZ�3v1v�j;�R�-��䘌�ܻ�.���T8�aݲ��-�,����
�W��3h�pě�r�%YyY����eNwu/��{������������!>؛%��ⴓ��ieVQױ*E.��w % ����Ty~�r_�VK��*�f�F�PXI�FUڞfjc��*��u�@`�o1&�O�� ㆊ/q�E��<���t�~�}p4�Y�{���'u��9�G���H�Q0ԁ(N��Z��FQ(  �j0+["3��i"~����ٌȎ.�6?���kdO8�f�W�J#E����[��p3�O��� �Y!�vȹ������(狙����Dd�
6]Ah��{�j�;�0(]�r<X\�uwʼ��#C�:j�d8�����5�Q�o��S�c��9iNP)�Tyt|_ɿJ�f��g�V�ڗ�Gs풛�o���l���B�M"�]��rX��"��
�$.C"\�N�T_�tf��7�@4C�'*[�`��ix���=n~�}6mw�M��cg}E�Ap
�`<�n��s�C�U;�U\��,�S!�7���l�~ꥑP��Q��p��=��{�X]�`�>�Ϣ{�e��u��:'���?#�%�F��`����0U��llӇ�Vb+Q,9ő�kX̄�F˥?2O�1�ԩ�폭j�B<s�QH
jK`�/�Ǭx�-������57k�[�ԮA�h�_��AԵuF��ƌ�$���T74'��[�-�d�Y(؁���\�/�T�2�$��f�Ot(�����k��ђF/g�C�Ƶ_r���!<��D熷;�ҕq<�؜C�(@͠�O:�RD	�5���7D�L/���iN�4G���`��i�`�̽��R��IJH���)Iz�+?i����� K;~�\��}M� F滔e~9d�O�Z2 zlzG=���V|35ħ�E��Xny�
����3X�aW/H��4��g�*:1LzS���8	��,ΟbK�W@���y�N"�����z��*�3^�v�}�N�-Ƽ��p��)�CD�W�Fw)�`��!�=�,S�5�� 	W������{��V�5�t�#?W�����%oͫ�_7�s?����%j��>#�мŉO5"V�?�֚�|_)��y�C�į�U��y��8'@�G�C�g���u~,1s/��S9�X��n�7 �j`aS����]�]�3I-����@�0N��YT.z��^ģ�[�����S�D�:�䏧��υֹ�0�sv����5t&}ބy+�Z}���:d���CH艺�E��ڬ���,��J+j������r�<��.���2;.U昈8��@��fe��%��2&L3P6E���Y.Y��묙^>Ū%��2��9w�]��ʐ`1�h�f�g���-�o&[ F�G`L�!��$Y��|Ld�W��m>Q���H�3�,3S�>�l ��l�{�i�C�I=(C�Q�]"{�$.`���j�}Dƚ�42��\(��lλK��6g^y�D1H�4ٌt�@�d��b�H�E�!Az顭KH1w�L��<>b(0p�Ϻ�P�����w&�(ҋp��>w�ݲ�Z*��g�0^�3�p������)��-�ӄ]L������}@��z)�����0���ˈx0�#����ض���� .O�8�;�Tj�!h.��xiE�aׂ���]`�G,�X<��6���(H5���^Γ]v��7��&�sd~k`wU8�(J���ǣ|�Q�9�����µR��h�Dؓ�+98�SʘÎ1]w�eIJhK����{?��wP�@�GP��!ДpR�4��<���|Cԙ�F�vr!�p&����Gg3�c�5
��5D`�I:F�YO�<��:�vbq�c�Hl�֍HF�`_k���[�n&t��r���O�#A�X���R�*����V%:�&��a{���2���_�̰RR�74}V�-t�aH��]MUBs�Jjt�}�#��9{�%b���$��mh徂F��:�^,:�?����q	<a�&߅[����w�x���n��@6�k��U��s\���1S!�{�r�!�����ZQ���419��T��G�y��4�&x}�L����w����P��`EZX�<��"6�Igx���p�Y�\t��$o^�E�D� ���I^\�/p�cǫ��8oxu��e�Jb'�[f4qA:q����ϼ�]W��z:�g�ܽ��q�H&O�B�z0�ӷ�K}�h-M%P��[J���Q91/��4��v��(�!�Ug���i�>���9�Q�]38wpwC���:S�F��8�����G[N�^��c.��.����.gn�3k��
`�*���y��I�=�w$|!0R6yK�d2���ah�؋�VX�jʌ��.u�U^���C�N�"gs ׁf����^�:���)<�H���`c5X~�bpzꔸ�-C*Sr���I���q>��ﲭA׃� �Ս���@�Eo3q���3*��:X�<72��qkJ�?ŞZ�w>ّ�^q�-;nĻ�(�"�q�ӷ��!,��3�{g&6\��
�x�Ӊ���􆌮��B]�3��-fA��/J0l���غk����կ�Ʃ|�6	R LM���f�i��V2F���o3��[�4��U�E�
���6���}xj/| ���q��%�`��B/�6�K��Kk6�8u���i�>Fʓh�8тz�m���W r6�8��>��x��&-�?\��cJ'�ݞ��ZY�[f����جGk*���0��@D�f�u��֮��[�Z#]R{�z㬯��S>���[B�p#S,��Xzy��ؠσ�9c��ARA��O��?s�5ᝈ�.���6'��{��(y��e'�����S]Q�w�l\����@3߭}9�@/�-�@���A��� ؔ�n������sD<��+E[�'��E$�lI���P'�H� ��
�$>�ld��9��da[wy]�G�-zМ�,�<��K�� �;�0Ks9��k��� �N-U�����C����u�����hB�Cʳ�5�w�(i� b4vjA��1I�=�7�jg���ݻ��WHA�<W����Jv�L;���l��./��ib��c�ޢ�R�I�����y]�H�ҟ{��tSXz��F��<�"о���yQ��B��	<��Ō���� ��~��t���$�w�VA����A mx��%)��e�c=��3�֧U�x����D]���Y ��`�:����G��ҁei���r0��B�LEA��7��2u��]���h�Su9�$���X^���x�QO��U�z���P�X𫂊�;�� �X����j��3��P��=��%~�iڜOQs`���o�i��Ǚ�XJ]���B��?�Z&th��VJ��
�\�|?�(���.w��Ȣc�����M{���瑿v�#��Z�U���e2�e�#Z�����e#˹��f���ND3k+�:<�i�v�i��Ozp~R}�((�2e��Z����18dFB�0i.�|�4����TZA�-��x%̦�o�C8UZ�Lʳֵ��^�L�����yJ��Gp���x�A���d.�x�P��z��}`�h�~Xl�f+�A.���8���4��>�v��!��|L
�e���z���,�Z��B�ِ����6w�=ﵥ�mV(놫1~�5�����n�I{'�/JV�i�?�L'�it��׼?�[,xUL�0 ӎ���k�������U{p>X��L-C�,[:�ƐL�x+R.�v�F�^��1A �ƶ��L4P��e�>��M3K��(�f�T�j���[M�1��5&!M@Qd��лc�J%"�� Zc���5�]=��5��P�I��#�x!d]��9�YW�"��=���ǻ<�ATL�[>����y��hq#��т<T����~�՛�=o��e+��*�`�7����wI�Ƌ֊i`�0�����@[�Ƌ�]��D��jZ�9��)�S�-����<�vrL Ȥ�x�+騂���|�w+>K��+�^�9mx�B���&>�L�'�U�ӭ{ng̗�-H����[�ʱ���+o��c`�����í��B>h�G���B�E��N���w(�}s�N4�!.��+�;3�"<~؁W9�;���*!�'���m��s@'�u.Ay|���JnJ��ƽ����O�$q .*��t��<�0��`�;�֚�r�1H+��|�5�@�'Ps�E'bGX5�����j:���@5�e|�qۢ:*N�F4�'ku]jƀ�3��J�5A����C�žE(��jgދ��L
w>�L~=!�o��r��Bk��rv�.(�Ƥ5����>��"�\k[)#�,^	��~���s���
\^���\z�T,6*0όD��z�hޒ\8ເ���rIH��&�G1��t��v��1"X�նX~{��;�����P�@�Kp��I���A�1�┠�a��I�����t�X�d+��^4G8^g~��d�4�e|��$�Ʌ��+�+�w�!K�<�ɨhf�%NyqW����׷�$y�G�Sc�T�_���3XQ�m��p}��/�g�ho|��B�c��~ڮ���\��6��/$O�y^�/��2��Hh��-ŷ|1`�,K�ұ*�m��m��w@���@n�q�V�q��~�9��>�X�»0�z��	��/�����_�>ia�U�9�ʞ��^>�l�@�j�1H���V-��|��<��� ���n��H[=p9�s�Ez0�y�h<�M)��ȝTeX��Yc"7��!�J	r�W-?� �:9D�,�����o �p����P�r1����2�RS���e��o�\:1wЙ\}P������ґ�o��Ө�e��8�'��`�tહ6��� �:|lN�'_+O.ri|~��$C�|�\UBy�Ǝ�����K*��m�4E??Z�Pb�pg�)c�T�C"���u �#�ov�^U�ϧ�}qS�i����Q�ȋ���F`:�p<*C^E8��k�a<(��uL�s��,�?�����q�c<"�ե������2D>�2����&�پ�m�j�H��8��ңۂ��B�&l�����L��9gE>U��#���%��1GY-ײ�6Y
���Z��Ը�z�Yw�{K������KP��lP�t��5��Uf��'Ӣn��^U޾�����=�ϰ����P�=����yU�F�w���A!Y�Ar뷻n� !�I�2i0�:�yA /ᔈ����e̪���R�� ���_��J�A���� ť��Ԙ����F���|w�|4M�!��|���2���}!f��Na~�ȧW�f}�<��-���V>�'#��g���~��E)�?�����g��;��C�,M��F΂Y=o�5E#��^�9R���,~���2���CeoliּwMN�V�W^�^"%��YD/�,N��K�����)��Q��]�ؼ8鯌G�a�u5��+ړ�R#ϗ�b{�~���<cV��F��	��-��j��[���p���� CB	�ۘ�6�`E���*�Z���
��4΍����8<y�����h��߄-M��F������E�u=��p���zH<�=�h����]��r���C�����st�'���8��0*��,���C*ѡ�R��Z�*�bWN� t�gT��u#ipiѲ��b���97AA�)Il��[Fg�$b��UoU/0�w�a�g�m� h�u[����Y<�����bd����'ԕ���a��
bk�F�-T6P׺�l�8�~�慹=�t({~2O���#w����Y�!���"�{���F���H��y;�d�LH댪w��ՊMo������;������=�K�'��<Ɛ��ߺA�dͶ�2�#��ŝ��20o��,�` MFm��R_�fg��v<!g�5���_#�:�����/\��Qh��ULj�̥�,�z������@�'�����`�#y}K�c�:�8���?��]N?X5�v�":B�~OPӀS��Ʈ'�ѡ��L������]�,v/,۾�_Ռ<ؤY�����{�������2�����>�GY.�f�Nj����.!r�E�A ��,���E�a��do����DY������^�_Z���������,8�i}�"ׂ����QM/³o�: �����\4�m!� l/M��^nſF����2��z��0�����V�����wE=�)��^�6QM��I@��_��pB��;�a��T�1&�L���ɃIg�37�z�t�_n`$�( 8��c�-�����w1�����'�Ty�������M��W�A�E.��Mt��t�-e.IxD�܉��w�
pt麃_�u/i ����sc8�����,1[qXq;%]�4���561�sȾ�dQ=��=����rG{]�wo`�o�c�,xɤ���dD.vZ�G�1wO"#l�s�gD���mU�t*p|C&�G��T�qt����m�8l�1��x�5ԣ2�o��b>�U�a0�0F�lq�_�:���t2=���T�b+���
�$��2������e�ģ4�jy��a8n�H/}��޿I��/Q��x�߃Bi.8:��o�:��'O���H�a�"K����r���&��j1�?>W����zo��MH�,�
!9:��Hݨ&&��~m�Tb�$��=B�c�/֑ß��G3�t� ���&?l11��M�6��S�W=?|��Y�8��Ge0�<To|H��y��KY6����l�S�5���hʀ�D]ʮ�{�=��m�W��F�>5	��	{ I�0i�.�����_W���b�aVU �R۰��\����}h�����x��$M�kQ�>,��%G5A�N��~��n�)'���@�H��j:�r�Ij)�Y��5�{��ܼ��PB��v9M�;�r���/$�W�mߥ,a�B����o['gxڹ������\f�	H"B�I�L �|
�ׄ<fM�CR�~!U]��I����72�G?.�0�3����P��8x�� '�`����� x�E5��䴵�;!)ж���W�I������C��O^�xs3���/��z�g&�Z�a|���)@���cu5�����?�֯~�\w:�qK!�eCV!���@6�lf�� �As���5Ʋ�q�GN�ZnD"߾��#���h��HT��@/�(#:c�v����*~���4����P�����Ë�-ܣ���}p�n
�a3��޲��"ӂp-������{�/��G�+Ph�}���b����1�h�w�C��-���1�����7Q�o<�:�1���mf05>W;��L���e<���l������G��k�	Ts��9���Ipv���4�}���*�]�D?��iLm�FV�w��l��3�c��y;�j�y�׺��F�
�sk��{��a��'�t��/]���Q���^�:�F,�ɊX�MfF���=�u���2$ ,������~~�q[�5��f��i��+1 �h�����^�`r�
P��`|����D�g�� d!@$����9��4r*���wLY��-w?�Z|N;�����ip��%#;�9��hl���ir�[Y����7���ddz�V�SB�j��ʼ�q�5I��^��=i��2�md���X��h\�!P���C�%	��i+f������h��D��9$�n4D��M�Br8u�n��3�E���N����Z�#�誨�T[�@c��y{nk�Bշλ��,���$]v�*��N}��I�t�|˲(�^	���kQ �H����ʗ1^ ���sPq%�{��;XP���u�|e��]��4���ɞZ%`P˟H���Ze)2#�	�a���4O�5+�r�j8���
U��ϻ�Z���V��q�DeoR������?(騁!b�R�G,�ܳ���'���R��j�2���H;X�Jݦ�J���Fܺ��z��ϿCW����Z�L;b���0F����Cy`[N����v��XI���.�-#7���w{te��2|0�!�c��:����ly�YHFH20?�'�Ծ.h���E��c[���s�Ĝ"�(�hF	O0��?H�$��c������,�M��L��ɲ����ьT|D2�ճ�Q&:Ia��u;�jjM�i�]{*�\�:��f�X�k!�Ü�x����R*�ߞ���s�����y��Kz<?x0�0�9�n�!�/�5l�"^3ɔD�7�T�Eoc���n�u�.QP:�lr ���)�ͷ���^G��QL|����W;���z�?��p�3�����+\�w�~��7�(n�"*���Uh��7���l��fe�����C�Qs"�=9�� �&qv�۲I	���$r8����dj>	��� ����1��Q�;�Hc�o�/l�rK1Ձ�=���0�G�������C��!hW��?c�DbE����fވ/v�^L(�p�EL	�l�^"�"<*�<�T^Ք-�*/���$M �����_���#j�-�w�
��\̺c�-L9��Ԃj��1�_s:̒c��s�Orw��\nS��t�!8B����e�*�L���' ����}��rP��j�10�OQ���瓃��o�n���P��`Q<5���r�������`4��y��-Rm�^rOC�� �]G	�YQY�BQ���d�rR��	�9@�C;F�~rk&R���ň��+�k��֮7�Uq��Qn�ֵ�'|��J3�o#�)�l��/�I��wz�*�t�e
���*S��J�z'��+"#N���!���>������'�G��\�Z���Z�㐙�ؗW6��F���!��K��|��o�~��7�.��~��H���v)\�҅�X1���g��6�+����Ra���2wi�����B
ܽ�N��etK8L�m�l�m��\:r��<j���Ѿ��� -�XS�;Uz�rJ�䭲F(y�d��P�,;?
��&9���0;Cѻ�|��L�����RKJQ�Gp;��Xz�z_b!�z΀m`HLN�Н�3����6��`���CB8ž'#�3H��A���Y��8�]��``��*^d��9]N,bńu����,�o�p�	�������8<|���R<��=w����Ԣ)N�U��/�/��ȳ�~p����6�]��R������%���p��7�Y�{v�nuW' �[�h������y�߆ߢ��P�G� �+�����1��ڢ_5���J�����/L`/� )#Ϧ�T�حޞ�I�����M�J8V�.�ۿ��W�R3��%e��Ž�`� {Qu���2�V�A�/��Y��$2�i�H/����BpcS|�\�N�+	�t/���e�/�4��$�����fH���2�����}�dV����B9�H^�ʇd� �<	��a��0I>�����A��h�JSw�*_��{���o�rKT[A[��-��="Y��^Ƿ	�jS,.
0�]~Rvi�9�m��j
�!��o���ɦ�âm�_#���ݍ.fH�a�!�
�tYçNՖ�
��87���IR��Z5PFX��6!ܤ߮I�Ar����ٍ.�0阅�s��X�K�B+���H8ˎ�j�vd�]��/f��Am�6�x�q�W���n�V�2������MN&
I�����Ћ	��zv��ef��01h��&cLH|;:u�U宮T?9�\�J(��M]��
�$�H:���엹� ����^c�0O��9H�-mˢrv��}ڸ�y��ڸ�E3�^���5qo�Cy09�4��n���Ǯ����4� I���- Ux�E���ӄ��F�y��3_Y�#�̝4������|���^��6^ɅԘw]���+��Zb��$uY�H�tq�^;����Bېھ8�v�ˮ}�,[3��5}�#�P���ۛ���D���k��|j�p͏$�sl���hu�,��t��&%��p��m�q�N�v���X}<Ps�_�iyWex�@�P��q�N�s7�
�l��Գn��=������djs�A�n����Fs j�W/�$���l��G��W�L��iY* -�M�������-_����T�܄q�q��4�c��Ԝ�lw#���|^�u��M�qLۦ� �DT�H�!�k�!�hRS�$zlm<vp�O�	� �્�YFc�~�H�D�|��L}�=AQ!��4�x�ɼd�m��@���N t��m�~��4J�Yi꥟�Zc�����y)8��̡1\H�1���{_��1�~7��x����É3�XB�Q�O�4�ڢD���&��g�2X�MIf�<���oq��B��\��OD�Յ5�ZΘ�y_t��ో]g�)��J���#�\Ү+k���$Q|A�잵{��:6i��Sť�3���o�<���.$�W��E�?��>�!OŃ0�@L�n!h\�%�dA�r"�2�d�>j&]��pB���2o��3���C3��AA2��/�Y��6��z׏��Ao	�����G1x�?6H �\������7s>�����p�c���CX4�����hD�2h�t�Bɞ�
��`�`:
{;k�yrT��jc�w�)���Nɜ/�Q��1A�WO�/�*�����ң(��f��5a��?BU-Xca]~��cy"Xk+�4�-�Z�n���F��n����q5��kd��D%>9����N�#P��յ�oHse7]��x������x�,�.���-��/Ӫ�B�}�y��ˑz��ڏ26S
�U�g��;9%ug8���VQ�$u�wv�Ym������6.Ơ-ӣ`�mI"�'�)��>��
��߷~3,5���ܥa,��f��Hj�ż�:?��S�m?w�8�l���~��Z̧��{���nZ���'�=� /Dmg��Pr��o�Q*WS�A�{����\�����b��mq򷒚�p��EU,�3gPp��T�\>�� �������8���a8�Z0/����cu]�jx�#��� ��$*T�Xry%��Otd���1��vah��l��m4��K��;�$s%����56�>��X2�3�y��sG�GL��1�y���������1���]��1�`�ǥ{�p���_{M��
�^܂��V ��c?Bf�^��$�=q�o��^b ��h�{,�l.� t�Dk�m����\�%^���`cS�x��f5�EJ1<<����t/-����)}g�	�P�tQ��'|��+X�b��ƭE lēm$э&�WH�xg
x>�ј*^Q�p�lU � �e��uDe���3 �̵�[�+�ٽ���&�{Oxw1J���=�+ҭ�43I���vM~>���^�3�v���=<�����eZ��tĿ��	�A>��.pʝ�ݵ�MG|�	�d�~�?�G$Ն�܆B�����%v��jB�t��9�I$�f���DL��!{U��C��bGg��^��88L�l����qa2NcbB�d|�%b_ U�sk����� ��=�`X؈�Y�Ӽ W#���M�ʬ��_�������_�ag�!]�8��6R�}��[&�AU͔�|� �	a��z,�{vf���1F��-V�A�
6A���}h�N�b0V�u(�Rݨ
o��2ᏨF�vC4g1�R[�e��^�����L���h�:/T� 5��"�Y����	'`\�d��;$e�4��%sj�̒�X�+I�E͔ޅ��\����ZčZL���k��ф� !컣ζ
��;�M��1B��f�5���}�(�$�]�H���� cK^���j��������:���a�C0	º+�f�ג>%�	HP����q�)�z����kb'�L��&�vxJ%(+��z�54]142��^�pM|��*���bh�+�.n�
w�|[���u����L��O�����cL����=�O���1F$(2 o��X(M�;�/�	T�����4}'y�*j�!��#�PEW��n���jo�騎�g K��~���5-}\�iEt�'��42�+���5���2�f����>�nҧ�/� 
Y1E�����r�@Ê�{��C�ԅ5�����;�G~���b��]��|ӳk��Ǆ������[�3:���%dJ��7;Xm-ܛR��'es��Z0w��T�'
l��D��/r�Q���))\���;�pҨ�~1�#»c�>|j���s��~��#0C�_v�5�2J��HȻ�≈�G�����/��l�-���c�j���+�	���ږa�}AhtltPj�`��k �Þ�5e�W�9F�G�����c���e�4��Ɖh�}!�,��o{����cL���s��Qd�bCnGS�`A��"0q�6�H���Fu�7bG�s�~�#@
3Lk�p�څ]K���*B���>8��'rEV"���>��HM9���B㜎j�<�4�c
~�.^��*Q�-� ¡^#X�v�̑w��3{���_۸1��>auC���:a��Ѭ��N-K}6� :Q�f���t���G�1��[<>6�o�g΢�,��*#�p��!������r�.��k�"�D�!��+�2o��~�R�����mu�8�3�w�pY��[�"�aK ���-$&5��˂��u���=�z.����2✷��]�:�М��řBb�� 	��*V8�ݾRQ�uR4��%��x��'��E�vO쓒���j��ZG���0^��I\U��eB��) ���~��Gr����4�$UJI���f;�7=|n9���ͧg�o=	�e2�WTr{�[Y�S^H������'���{�è�Pp$�;�܌��@?�7BJrm��L��#�E�8��/�3
�v�%�o˽�\�f�e�T�𥂼4:�^���jR#]�38f��@歆���z�y��-���@ZC';����J����6`�[Q?�H{�<&m�����jg&M'����l�3��R��Y��$~���?�t�q=��~�'��û)�G�CD�2K�S�_�\fop��V��[;~Hh˓�m瀳}�CE�;�4ц�=�7_g1��]��o��Jq H��&
���Y���xQj�[�5��~W�8�y���v��ߑ<��bt"��=�bJ�˽說��貔�M�k��-�׏;�F.�p}�֪�	d����+�9�v:�&	a�ۦ�l�U��K����/^Y��,v�OIX�T<�gs݌��I��Gyt]�{ӳf��ǵkqC��N�0M}�7hS݉��$�u�9t'Lu���[�� ���-rPD-吿U����0Z�B�^��NW��2"v]߰B�|�� ���jz������pL����b�c� ���o�/��ρ4?��@lP�?�����?��i[{�<R�P�}�z�lϙ��2 ���|L�*���T�B�����c-���q�v�\O΍��I�.PS��hʟMBZ�d(7!����~,�
X�
!�${��`6�>^�KB9���j���6��Qyo��|�ST�*Y%��&=���Ǫ:����w}w�G��Fɮ��m�PKݵC��y���j"G��ñ$'�S7`�~�۰Sa� -7�b+9��5l}6N{K��c>�%E��"�?4jbl�5ZN"�����Y7�d�ia#��!�p�k�Q�;2Y�>P�o8��.���[q�Q��6-��KEq6��YEx�Xj�9fA+��V���8|�M�b�L]�����F����j��Z����L�U~�Z��.!�2���b�o���Id�7�VRE�0� �V�Z�i5�,�HW��X^�P���v�VP#+q{��,��Ad��.5z��ݒ�=o��Y�[�#��R���y�C�nK��b����q���ǿ@��:�=�����0D���w��HGkbi#m܀���38��f99�.�Ν�z�;���5��"�,<F��.��g��e;�5��
<(��O�JOe�U4H�;�'	�.����Ob�'r)8AC�H!�R�h:"�c�K��]i1`�S9��=Ɩ���gI��ک��4���m>ᴏ2��h�9u"u�6I൓/s�� ����x��/8�0E��DN\�<�Ľ���94jn~��������{�MR&
�)7�j�t�������f:+9G�;_9�����.��4Gƶ��3�5�	T���LLO��Tw�r�CAK����el�N1���Y�QRq+�qvYm,���Sp@���8P�RqX�ac�2��Fz5Qg�����$��W�'n��e�9�2��n2b�VI���]Q6��-�r�cF<�)�rDZx~kϮ*[4��{Θ�]A�QD�����K��Y�<-�*��1�1�\��
�R<�^�-I^�hj1�Ź{��:�m(x�A����K]�X}mtl6��;��i
������a����Ny 6�Mu�a}�c�j&�!�cK���7g�����?��T����ׄ<����=�Ĵ��N��^�K����k�},�@`�E��������� �r�K/.9*h�-���ĻbH���<`[*�vDKQ�F6�|�|�hTP�׹T#�5����!��[H"(1�A�]��61N�%A�-��q�d�!|�^�dp�W�&u@�0CW ��įS�K�f���|��J$�b;���e�F�>����m�#��O+�J��yi?	��w�kO���G��h��du8dl���?M |��I��΁��3&�ԚU�}#�{"�g�z���i�3�z�e��%�B�Τ��Dx�2��	��k��&G[C����"�w����͵�;ތk��ٴ<ʤ�`m;��SB>�}�H�v+{'U�����=��>*�pQ��
L�^�α:��Ŭ�i,��*�x��r|ܕљ�����h��Uwܝ~ �08�
D0?Vtr��a�R	c�U�,@�J�������0�Y��,��#!�ʒ����O{�e�H��Xb*:��~�+��۸�#J��0 �aMF1���&4��/Q��2S�m�p����5g��ܵ/��	��@��zqM��C�Յ�NF>*�;�����Y�C_=��>n�<�y�4*��p>��c2"� ���Knb7�9�Z�XU���9�`�)��eg�$��1����I�M�Џ�\���Fҏ�8~|O+��$x&=�ER�iLM��N����`�Hf�O�x��>8�:%��u�m/U
�Hmhz��+�9b]�_Y�M,��s���@��X�W_���F�6r�"��������DQ/P�9e��L+��)��r垗�J�`�8{�Jf�N���hl�0�0�n����I�3ep��;ѹ�;�T�K�M�~�R"��*��&p9 �
T��;9�?��~���ϽV$�3z;�7s���NO�6�wt��3�PF@�uh�彋�I��΁�ԇ0���&�q���N�O_��:x����T3�bU!���y��cFo�\�zG���w����o� !'*��}�|�#�-I%}\~R^��B��V�_[���k*V�>��DlD��8=�K RW;xJP)��o�����=k�ں��3ȎMGGL�����{���{���pk�Yd�&�k^0��k��q��ze_r���SB��t+w5CC���͌�����-�Fu^t@!��*�L��l�Ԥ��9��ig.�,R�3�f�r�]�3���%,t��~^>s�?�Ю&b74գ)Zf��^E���5!yR#��v�� r1s�3���/g�}h�;N��^�D�*x���Uc��V�ML�>Sb/�bV�"�v�ʿ���� Ak��ʠW�����U���[���@3��"���=��tF���� &���*�n�����Nu����N#kQO�3�ǹz�a�o 2�Q�������doN	M�Qً]�q<(�2�e���;��2���2�����URx7����BB]g�����9z��N�`h|�dkͽ�ڮ����|>�/�`��c����wRU�O��[6��*|�z�ȫ���NR������������lY���l_K��]�l�,D�\�'�"Ndj��������h��2�0M]� pԨܝL�q��o҈��4�f�f��U���(��M�:�Sl;�����.�ŧHV�����ݻ�=�=x�O��e}A���dwu;�Z�?xXfnF�h�	�C�Jq��E`oޒ»|!��z+;˱`��c���M�,�o*���>FL����DIT(��7���j��i�c[=�Y�*?U=8`�]�`²ǚ'��<��9ɿ[, �C4x~/�:3���U��љ�~�EN���У�i<����*�4��5��I4|��2+&���i������r��W��n�|H��K�]�ؘ��^Qm���,J)�֊���H��I�T��������!�\U���w��^8�#�1;�h"�m/I�ɲb���p� [N�@���G�>��!�|cg��w�	�����u
����°,H?��̓�7K�P�:v��W������I. ���"���b�6��Ý�{q��AQ��&a�Z(���D�;��[���A�=�.nC2�CeVy���E3��b���J�G����!ҢA3�ЪY���'�ق[nd�R��5��8�,��PTPY�ErZ�ݍ���^�e�K�������B`��BH�A��y�������竃�}��w��a7�|_l;�yF�A��B��H�"���+��u\Y@ép��#���X�6R���7���2��O%Pu��j=Y/�\�k�t�:۷Ӛ2�e��������G����N����tiW@;ʀz��a@�a�{��=���Z�Yh2�`*�ÜИ݈s�(u���H��{1�	L{/����0����/So9;���a
�(�d��Qh#�R�~�c!�q4c�~ц?D+aR!���#gK{%��+¿13��|d@������x|��[-���a�2�}���ʍ]h�����{m]�5�ǈ�jC���^�`y�$J\�v��j�4�iw6���ƞ�Yl2OGF������B�Z"�*՟.ii�0v݃��e#�[v���F����䐊 ��Y�VvL׵y�� 䮺}��=��^2UO#>�?M�F5��2}x|�@ �A��	����	8�����@��0�x"�Oe����x�7Uը�B�^~V��|(�h����-|+�#O)�P�FcsʁZ  ��-ՔF�T5߆�7db�En|Qz6Y���«.�6DdgD����"m����!6��� ��	��^kw��.�%7U�F��y�df���(rG��n��Hf]щX�]�RW��#�>��)�ybI<���pI뇤�q@����8&��>�����?H�L����lX��ݖ���T�U�g�C_Q���ű<Do�|��Wy�ޫ�Q��ؤ>U��D��4&h[փl�t��xP��s�~�,����7=?�?�?(6�O�ԩ�I�7�0�O&0=�X"q�������
�[J�uΑ�<���A��.��T�j�ŏ@Hh�x�����ͣV�����e)�g���)��b��Pz�|R��j<���tL�����w���N�\f�OL�j«M0Tb�El��5a��2@�j��F�9Ɵ�->��y�7�nL����r���)�Vt'��p�i��{[Pi���|�����u��?�C}��)[�X[��1������˰�wSP��6��6͡�8����H��I~��8ĘB����H,!1��`Л*�i��e��?�!ư�,���і?���*脭�����;ʔҗ�ǖ�\d�����[�;��k�E)�嶇�M�J���)Ԇ�iz��
���'5�'�g�M>���qf����q���O̵���;l���ב�.�)�D\��w?������b5�I�h���T����D���V-�!���
�1���FQ<�ln�n��F�����;���Xx��:�7���_��z�ٷ��&hrp�f����\�*�e�O��oX������( ��^��<��+ $pJ˝Y2WJ��\d��eh��W�w��Ҍ�S������ݛŠ��4p 2]]|��q�jc�1R@F;W�u�'DSa%fT�;�}^�Q���V��OO�bO���}�w�H������}p6T���r�ME��y���@n�uO�恎W�x@9ĊFּT���e���������t�w�I��H'5Q���*cL�5Ta��*F@Q�e"�R��9���(0�)=��X|+=o>�hB1�q�a��66T:�-ؙ迳�f51!hr��Ul�m�H�
�R.�=�=�}U>.�,v�N�y���Q�,�O�y/޴k3�y<֟]�s@,�ҵc�ߏ����Q�"P�$�����,�&���Q���F� ��߽ۘ�[&�(��o��-�(@��8'5���,�]�(���9�N���j<����8�D#qP؋�zyip0��ƣ���#��{�x���NV-�s��$��l��j$#h@5u�`�6��Q�q6������e�ˀ�U�
�3~_X� ��H
K��S����vX|������G��/�7������&N���S����x����7{���M9����=AC�0᧴2���h)�M��1��X,��b��b�{�pZ�#��DʞU�����d�pip�hĠ��朜�݊�h%Iz��6�-�`�6�+�F�oj<��31������g�< %(-�a7�!����x�p�aybŕ\(6�ݫ��*.����pN`j�h�t-�g���Үt��})#���@�GIl�\/��?�ŚȮ��/`IZ���<���V
��ľMM߼֌ɥ�|J��ݔf��(Sp�ݦY��{�ބ�=i��
q���|����'%�?�u#��*@���RAuހם$���xV%�xU�[o�*�G�B^+q�dqf�-f5i��G�i/�(`[��|pX\k�i+��:9�Tp(�V�d��ע܈���^(�G
o���K��x�cd���.sAnUA:�(t�)�4�&�<ufY���M�=���ش3*���M�� u���ǜv)_.����:��_X`K{L��K%\پ2��q��V�7i�36��R�-ϸ(G�sVY��J�I��΍D�޵�+��F������  _*f���.���=O	�¢��u<x@�0�UDh�*�5/-����,�G=��)"�;��xwjs�8?��h��CА
ِ�-Nga��u���`���4���^"f�?�,�s���Zk_���?��p���������)lI��XT��1�t	����j#º|�zuÈ���ZN��V�_@ �aE9->�mPt�=�^=�S��h=��!���7xܦ��-�t�E<
�?���D�(W���?�^��u��޿��UV�z��N��FX�is��Y��O��O���X�=�u�p�)`��̞%����F O249��=�|XF�����_ůy�aJ'��`����"{�u��w� ֟��y{;(�\R�m��"�i�[R����h5�(�ix&G��FL�!$�V�Qʆ#h�a���U�o��b<z^o3�C�yo@
���,k�Y۠�-墓t�ey��hL�<�Z�"��#SUBI�;�O�[���h����fJ���˭r�����I�T K5���:�g�?�������G�,��Z��f�: ��*�ҳ*�9�T�9�%<n����n���v�~�Lyy�=_�<��ް�C~���hX�В=�uw����=M[�D�uu�t��6���9�8��Z�O�~�J*5���WU�3��s�j��Ҍ��6�=HhS�Lь����b4�L��u��S���*��W����-Ai�r����՟��b��v-��D1��!�.q3��0.yz����]���B��3!��[q>��Iq�d�g5��'�
��R�i�K�?U�1K��RM]��UA��H1�b�w���?L��6��Ϩ/`J�[Җ����ɕzS��m�4/�K O��!���P{b�i>M��Qm�/s��H�	�(uR�O}�� �>>!c��	��Ǳ�>/@k�+?�sq~�G%�������2.0�"ѝ�cz���1z|����^9�Ҏ���]z{*c�=�jt��?*V&]X�ܝ_go'����K��I����ˇ(+.{OvSd�i�4o?�:��}Jv���h� �%kF�d�qh�Q7/��r�����!��aN�&]{��q�%�~�����2�׏����U�-.��u���{)��|��z/��Zk�T�t���ZP5�1�}�^�2�)��k���^?�{�+&��")BU�.B�  �c%�M�ҭC�h�&=�jW*��	r����ӽ�?�o��Ե`m��M�Rl���Qe���{�6���M����#��>1����-��$�Z�Xs��TSbS��8$$J"�N�1�o������pbOq�"Q��$I}x)�qM%?��2pl����9*��ʌ���b�#�{~������q�"���)�P�0U%§��|KN��V	�~�ORr��e<c��y�"����c`Z~�'|G_ra��΃]������A)�b�}is�[ q��� � :�naoYc�?�i�`����u�&Q�	��PNXj��e&qY��p=ujW�S>�*��c_�o��X*5t��s����12>s ��$�ɼ�%�\�y*�)|!�W�}GS�g�d%�cC+n܁�Cm=�&
�#R7/EPI]�g4<��ܷ{5e�zE9Y��x�1�B�\pA��n�f48{�,���, ��Z��#�2F�c�9��z$ؼx�y��@�p�-�i�4�
���.P1H��nuבj����"��$�	'���-D^�xRk$U��^�f�S�V 7"�hH�(�,k���LmY�)Be��PH��Y]Aط�.x\L'�/���t�RW���]=\�tYP�D��f՗�xV�_ġ}�l��8�ِ�B�O�Ku���Z��`��$d���3`�$�U����;�Z��+ "�i�w��Jiٹ�IJ<�,���'� ۋ Ѐ�l��ܫ�o�ק�-�O�2��l%|`k�$4-�j�W�Μ�?w>�����qB��<�|�ָ���Z�00��3.��.�"¤ڦ�����W^�F���������d�ޝ�D�NG��ؖ��`�)�Y�RC�Q����v-?d
URE�_�o^�㌍��*Yz;�2�,g�rhp\-Z���r��Ҝ�0�H���|�R<�T.>�����O��d�߅(�K�J�A��/C���Oqti��Ͼ�E)���T�Suu*Z�̿�gVK$v2�����%�%5h�'�4�b&�:ȺE<��?�SS��t�z������qk�Xշ�~=W`�nE�i�UAZ��~$@c�	�]?f�c�I,^<���-c����Ό�v#4D���UK��U��R�5�rwdwNG�7s�\��G�(C�u�p��ew�PQ�i4\C��c�3���B���үŎ����d�WV��P��y�z�y�TaK�(�#Z��cX 4\�>�hUƚ�QQ�RИP�-~�7l��K�	�\�ृ�u*�첑�u�x�v�E�%�'�D�-8�4�p�ʟ� ."޿��P���� .�L�9�Y]Q�[wn�I�@�"���h�� �w�G;f���}�
���~�xc�₼z�]���^�c�a�~��oѦ�k1�إo�G\c���î���!�H�M�*�N�r�m�n����O.��^EL=��@�&w#��P\Y�n��;eѷ�wK͌:R.YF�+6�OP��Y���CZ,��D�r��b�Ĭ7A-~�퇧<N|��R�������v�Sln�(�� �/cE����?U����h��3y��!��?\�W�~�����?T�Ɛ�á�'�|�&+.mL
>�J/=>�Zg�d����\�"/��՗�v\��Ӌ�q��0��T�A�����wk�a=bzX�xHt�^{�D��l���S��3d��s���	�<�=V�� l]W;V����k�K�\o*��,�%�M��/6$�Ƿ�+�������06J ���L��%d�v�F�`ڦ������Q=Q��3�^����s�1=�I��j�k}��U�*Y^�_��	��*�y#�7�z�C�7P�x8N����rL�!�i�M`L_������ �B��w���Fʱ��A�i[��t��eo�tc�ȵL�[�jy���f�+���?�U��e�Q����[�sL �����Yb���##ƙRR/R�y�d����3��A���Ҙ���������-a�(��@���-Nt��"���`�eP3���t��+͜��to/���]e���_[��?~)%��W�f>Z�l(���@D�΋M��0u��GXgޤ��5�2{Bz��ۭ'�h�]Ot;�D�����9:�B�h�O&�)�R�0���[8�nC��k�۶�m�����
Z�(��_!�u�u�T���mPs}�[T�"���m01�[�uLĖP��~�1!(��'�(�_Ǯ[�Ͱ�ҝ?�1C���g�_1�	���6�!wz�Af>���=���D4mI����Ģ�/��(,xn=����`n����L��3���!G��w�7O�Է,����}�Q��,�ΐ��E���]l_���A'+�(���z/�T�T|��l4�*�ڪ`�#R�r�=�6]�V�=�&"�W��E>B��P/<eߜe�^0y7k�����{cd�q��&�	$�*P��O�,:E�o!����u������jFw���gt�$@����E�~U�U��U�P^��G)� �*�`�@��=���|腀V-����c����ș��8G�Ș�;�����#�=�a!�k���-ѳ�l?�����9��g�Ԓ+�?#�m���`5�4
oT��+L�O����e��L[�F��U�<=��ҝ��5	���)��'���v�
f^�yۗ`�^`\����y�DD9=��(�y�DB�_���86U<����f�
.6�	�j�6���f�.�?���vr-C�Sx�1�8�"�w���5}YL��|ۊ�)gr!�*��ǃ˯O=v��f����7,Hj-,7勫��9@L�����@��:�ST�K��ň�%)zr�d+t9\)(n;7���$?^��]x^������-VƓ���he�z+x��7���Gp?���w�N2u�g��6u,Idn���J��W���7�b�v}�`$j��`?*�� �V��94
<N �w(�ջ��'B��ߺ]�D$>�vjAh��:�
�N�Nf)��lB��s|�ň��" y�1.��hJ�E���ͳ%{�H��� +t�L�Ko�i�Hl�g�WC�S�;ZK3x�[��,�Iv�ٸ{B���$�rlx�ӿK�B�w�Ls�s�!�&�a<�QٕW�<`*cz���%x&6f�qL=��!��;���$�t�l�[xE��"��6Z&̂k@���wqd{Կ��vF����a� �#���$��2�ϊ�~E"�)Q��sJ����d
�覬N��3�����,���9��QC��:�-�,a�Mt߫��% D�m�p���p�x��;RmX1& ]�	�